

module test
(

);

  reg CLK;
  reg RESETN;
  wire irq;
  wire [32-1:0] maxi_awaddr;
  wire [8-1:0] maxi_awlen;
  wire [3-1:0] maxi_awsize;
  wire [2-1:0] maxi_awburst;
  wire [1-1:0] maxi_awlock;
  wire [4-1:0] maxi_awcache;
  wire [3-1:0] maxi_awprot;
  wire [4-1:0] maxi_awqos;
  wire [2-1:0] maxi_awuser;
  wire maxi_awvalid;
  reg maxi_awready;
  wire [32-1:0] maxi_wdata;
  wire [4-1:0] maxi_wstrb;
  wire maxi_wlast;
  wire maxi_wvalid;
  reg maxi_wready;
  reg [2-1:0] maxi_bresp;
  reg maxi_bvalid;
  wire maxi_bready;
  wire [32-1:0] maxi_araddr;
  wire [8-1:0] maxi_arlen;
  wire [3-1:0] maxi_arsize;
  wire [2-1:0] maxi_arburst;
  wire [1-1:0] maxi_arlock;
  wire [4-1:0] maxi_arcache;
  wire [3-1:0] maxi_arprot;
  wire [4-1:0] maxi_arqos;
  wire [2-1:0] maxi_aruser;
  wire maxi_arvalid;
  reg maxi_arready;
  reg [32-1:0] maxi_rdata;
  reg [2-1:0] maxi_rresp;
  reg maxi_rlast;
  reg maxi_rvalid;
  wire maxi_rready;
  reg [32-1:0] saxi_awaddr;
  reg [4-1:0] saxi_awcache;
  reg [3-1:0] saxi_awprot;
  reg saxi_awvalid;
  wire saxi_awready;
  reg [32-1:0] saxi_wdata;
  reg [4-1:0] saxi_wstrb;
  reg saxi_wvalid;
  wire saxi_wready;
  wire [2-1:0] saxi_bresp;
  wire saxi_bvalid;
  reg saxi_bready;
  reg [32-1:0] saxi_araddr;
  reg [4-1:0] saxi_arcache;
  reg [3-1:0] saxi_arprot;
  reg saxi_arvalid;
  wire saxi_arready;
  wire [32-1:0] saxi_rdata;
  wire [2-1:0] saxi_rresp;
  wire saxi_rvalid;
  reg saxi_rready;
  wire RST;
  assign RST = !RESETN;
  reg [32-1:0] th_ctrl;
  localparam th_ctrl_init = 0;

  complexcnn
  uut
  (
    .CLK(CLK),
    .RESETN(RESETN),
    .irq(irq),
    .maxi_awaddr(maxi_awaddr),
    .maxi_awlen(maxi_awlen),
    .maxi_awsize(maxi_awsize),
    .maxi_awburst(maxi_awburst),
    .maxi_awlock(maxi_awlock),
    .maxi_awcache(maxi_awcache),
    .maxi_awprot(maxi_awprot),
    .maxi_awqos(maxi_awqos),
    .maxi_awuser(maxi_awuser),
    .maxi_awvalid(maxi_awvalid),
    .maxi_awready(maxi_awready),
    .maxi_wdata(maxi_wdata),
    .maxi_wstrb(maxi_wstrb),
    .maxi_wlast(maxi_wlast),
    .maxi_wvalid(maxi_wvalid),
    .maxi_wready(maxi_wready),
    .maxi_bresp(maxi_bresp),
    .maxi_bvalid(maxi_bvalid),
    .maxi_bready(maxi_bready),
    .maxi_araddr(maxi_araddr),
    .maxi_arlen(maxi_arlen),
    .maxi_arsize(maxi_arsize),
    .maxi_arburst(maxi_arburst),
    .maxi_arlock(maxi_arlock),
    .maxi_arcache(maxi_arcache),
    .maxi_arprot(maxi_arprot),
    .maxi_arqos(maxi_arqos),
    .maxi_aruser(maxi_aruser),
    .maxi_arvalid(maxi_arvalid),
    .maxi_arready(maxi_arready),
    .maxi_rdata(maxi_rdata),
    .maxi_rresp(maxi_rresp),
    .maxi_rlast(maxi_rlast),
    .maxi_rvalid(maxi_rvalid),
    .maxi_rready(maxi_rready),
    .saxi_awaddr(saxi_awaddr),
    .saxi_awcache(saxi_awcache),
    .saxi_awprot(saxi_awprot),
    .saxi_awvalid(saxi_awvalid),
    .saxi_awready(saxi_awready),
    .saxi_wdata(saxi_wdata),
    .saxi_wstrb(saxi_wstrb),
    .saxi_wvalid(saxi_wvalid),
    .saxi_wready(saxi_wready),
    .saxi_bresp(saxi_bresp),
    .saxi_bvalid(saxi_bvalid),
    .saxi_bready(saxi_bready),
    .saxi_araddr(saxi_araddr),
    .saxi_arcache(saxi_arcache),
    .saxi_arprot(saxi_arprot),
    .saxi_arvalid(saxi_arvalid),
    .saxi_arready(saxi_arready),
    .saxi_rdata(saxi_rdata),
    .saxi_rresp(saxi_rresp),
    .saxi_rvalid(saxi_rvalid),
    .saxi_rready(saxi_rready)
  );

  localparam th_ctrl_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      th_ctrl <= th_ctrl_init;
    end else begin
      case(th_ctrl)
        th_ctrl_init: begin
          th_ctrl <= th_ctrl_1;
        end
      endcase
    end
  end


endmodule



module complexcnn
(
  input CLK,
  input RESETN,
  output reg irq,
  output reg [32-1:0] maxi_awaddr,
  output reg [8-1:0] maxi_awlen,
  output [3-1:0] maxi_awsize,
  output [2-1:0] maxi_awburst,
  output [1-1:0] maxi_awlock,
  output [4-1:0] maxi_awcache,
  output [3-1:0] maxi_awprot,
  output [4-1:0] maxi_awqos,
  output [2-1:0] maxi_awuser,
  output reg maxi_awvalid,
  input maxi_awready,
  output [32-1:0] maxi_wdata,
  output [4-1:0] maxi_wstrb,
  output maxi_wlast,
  output maxi_wvalid,
  input maxi_wready,
  input [2-1:0] maxi_bresp,
  input maxi_bvalid,
  output maxi_bready,
  output reg [32-1:0] maxi_araddr,
  output reg [8-1:0] maxi_arlen,
  output [3-1:0] maxi_arsize,
  output [2-1:0] maxi_arburst,
  output [1-1:0] maxi_arlock,
  output [4-1:0] maxi_arcache,
  output [3-1:0] maxi_arprot,
  output [4-1:0] maxi_arqos,
  output [2-1:0] maxi_aruser,
  output reg maxi_arvalid,
  input maxi_arready,
  input [32-1:0] maxi_rdata,
  input [2-1:0] maxi_rresp,
  input maxi_rlast,
  input maxi_rvalid,
  output maxi_rready,
  input [32-1:0] saxi_awaddr,
  input [4-1:0] saxi_awcache,
  input [3-1:0] saxi_awprot,
  input saxi_awvalid,
  output saxi_awready,
  input [32-1:0] saxi_wdata,
  input [4-1:0] saxi_wstrb,
  input saxi_wvalid,
  output saxi_wready,
  output [2-1:0] saxi_bresp,
  output reg saxi_bvalid,
  input saxi_bready,
  input [32-1:0] saxi_araddr,
  input [4-1:0] saxi_arcache,
  input [3-1:0] saxi_arprot,
  input saxi_arvalid,
  output saxi_arready,
  output reg [32-1:0] saxi_rdata,
  output [2-1:0] saxi_rresp,
  output reg saxi_rvalid,
  input saxi_rready
);

  wire RESETN_inv;
  assign RESETN_inv = !RESETN;
  wire RESETN_inv_buf;
  reg _RESETN_inv_1;
  reg _RESETN_inv_2;
  assign RESETN_inv_buf = _RESETN_inv_2;
  assign maxi_awsize = 2;
  assign maxi_awburst = 1;
  assign maxi_awlock = 0;
  assign maxi_awcache = 3;
  assign maxi_awprot = 0;
  assign maxi_awqos = 0;
  assign maxi_awuser = 0;
  reg [32-1:0] _maxi_wdata_sb_0;
  reg [4-1:0] _maxi_wstrb_sb_0;
  reg _maxi_wlast_sb_0;
  reg _maxi_wvalid_sb_0;
  wire _maxi_wready_sb_0;
  wire _sb_maxi_writedata_s_value_0;
  assign _sb_maxi_writedata_s_value_0 = _maxi_wlast_sb_0;
  wire [4-1:0] _sb_maxi_writedata_s_value_1;
  assign _sb_maxi_writedata_s_value_1 = _maxi_wstrb_sb_0;
  wire [32-1:0] _sb_maxi_writedata_s_value_2;
  assign _sb_maxi_writedata_s_value_2 = _maxi_wdata_sb_0;
  wire [37-1:0] _sb_maxi_writedata_s_data_3;
  assign _sb_maxi_writedata_s_data_3 = { _sb_maxi_writedata_s_value_0, _sb_maxi_writedata_s_value_1, _sb_maxi_writedata_s_value_2 };
  wire _sb_maxi_writedata_s_valid_4;
  assign _sb_maxi_writedata_s_valid_4 = _maxi_wvalid_sb_0;
  wire _sb_maxi_writedata_m_ready_5;
  assign _sb_maxi_writedata_m_ready_5 = maxi_wready;
  reg [37-1:0] _sb_maxi_writedata_data_6;
  reg _sb_maxi_writedata_valid_7;
  wire _sb_maxi_writedata_ready_8;
  reg [37-1:0] _sb_maxi_writedata_tmp_data_9;
  reg _sb_maxi_writedata_tmp_valid_10;
  wire [37-1:0] _sb_maxi_writedata_next_data_11;
  wire _sb_maxi_writedata_next_valid_12;
  assign _sb_maxi_writedata_ready_8 = !_sb_maxi_writedata_tmp_valid_10;
  assign _sb_maxi_writedata_next_data_11 = (_sb_maxi_writedata_tmp_valid_10)? _sb_maxi_writedata_tmp_data_9 : _sb_maxi_writedata_s_data_3;
  assign _sb_maxi_writedata_next_valid_12 = _sb_maxi_writedata_tmp_valid_10 || _sb_maxi_writedata_s_valid_4;
  wire _sb_maxi_writedata_m_value_13;
  assign _sb_maxi_writedata_m_value_13 = _sb_maxi_writedata_data_6[36:36];
  wire [4-1:0] _sb_maxi_writedata_m_value_14;
  assign _sb_maxi_writedata_m_value_14 = _sb_maxi_writedata_data_6[35:32];
  wire [32-1:0] _sb_maxi_writedata_m_value_15;
  assign _sb_maxi_writedata_m_value_15 = _sb_maxi_writedata_data_6[31:0];
  assign _maxi_wready_sb_0 = _sb_maxi_writedata_ready_8;
  assign maxi_wdata = _sb_maxi_writedata_m_value_15;
  assign maxi_wstrb = _sb_maxi_writedata_m_value_14;
  assign maxi_wlast = _sb_maxi_writedata_m_value_13;
  assign maxi_wvalid = _sb_maxi_writedata_valid_7;
  assign maxi_bready = 1;
  assign maxi_arsize = 2;
  assign maxi_arburst = 1;
  assign maxi_arlock = 0;
  assign maxi_arcache = 3;
  assign maxi_arprot = 0;
  assign maxi_arqos = 0;
  assign maxi_aruser = 0;
  wire [32-1:0] _maxi_rdata_sb_0;
  wire _maxi_rlast_sb_0;
  wire _maxi_rvalid_sb_0;
  wire _maxi_rready_sb_0;
  wire _sb_maxi_readdata_s_value_16;
  assign _sb_maxi_readdata_s_value_16 = maxi_rlast;
  wire [32-1:0] _sb_maxi_readdata_s_value_17;
  assign _sb_maxi_readdata_s_value_17 = maxi_rdata;
  wire [33-1:0] _sb_maxi_readdata_s_data_18;
  assign _sb_maxi_readdata_s_data_18 = { _sb_maxi_readdata_s_value_16, _sb_maxi_readdata_s_value_17 };
  wire _sb_maxi_readdata_s_valid_19;
  assign _sb_maxi_readdata_s_valid_19 = maxi_rvalid;
  wire _sb_maxi_readdata_m_ready_20;
  assign _sb_maxi_readdata_m_ready_20 = _maxi_rready_sb_0;
  reg [33-1:0] _sb_maxi_readdata_data_21;
  reg _sb_maxi_readdata_valid_22;
  wire _sb_maxi_readdata_ready_23;
  reg [33-1:0] _sb_maxi_readdata_tmp_data_24;
  reg _sb_maxi_readdata_tmp_valid_25;
  wire [33-1:0] _sb_maxi_readdata_next_data_26;
  wire _sb_maxi_readdata_next_valid_27;
  assign _sb_maxi_readdata_ready_23 = !_sb_maxi_readdata_tmp_valid_25;
  assign _sb_maxi_readdata_next_data_26 = (_sb_maxi_readdata_tmp_valid_25)? _sb_maxi_readdata_tmp_data_24 : _sb_maxi_readdata_s_data_18;
  assign _sb_maxi_readdata_next_valid_27 = _sb_maxi_readdata_tmp_valid_25 || _sb_maxi_readdata_s_valid_19;
  wire _sb_maxi_readdata_m_value_28;
  assign _sb_maxi_readdata_m_value_28 = _sb_maxi_readdata_data_21[32:32];
  wire [32-1:0] _sb_maxi_readdata_m_value_29;
  assign _sb_maxi_readdata_m_value_29 = _sb_maxi_readdata_data_21[31:0];
  assign _maxi_rdata_sb_0 = _sb_maxi_readdata_m_value_29;
  assign _maxi_rlast_sb_0 = _sb_maxi_readdata_m_value_28;
  assign _maxi_rvalid_sb_0 = _sb_maxi_readdata_valid_22;
  assign maxi_rready = _sb_maxi_readdata_ready_23;
  reg [3-1:0] _maxi_outstanding_wcount;
  wire _maxi_has_outstanding_write;
  assign _maxi_has_outstanding_write = (_maxi_outstanding_wcount > 0) || maxi_awvalid;
  reg _maxi_read_start;
  reg [8-1:0] _maxi_read_op_sel;
  reg [32-1:0] _maxi_read_global_addr;
  reg [33-1:0] _maxi_read_global_size;
  reg [32-1:0] _maxi_read_local_addr;
  reg [32-1:0] _maxi_read_local_stride;
  reg [33-1:0] _maxi_read_local_size;
  reg [32-1:0] _maxi_read_local_blocksize;
  wire _maxi_read_req_fifo_enq;
  wire [137-1:0] _maxi_read_req_fifo_wdata;
  wire _maxi_read_req_fifo_full;
  wire _maxi_read_req_fifo_almost_full;
  wire _maxi_read_req_fifo_deq;
  wire [137-1:0] _maxi_read_req_fifo_rdata;
  wire _maxi_read_req_fifo_empty;
  wire _maxi_read_req_fifo_almost_empty;

  _maxi_read_req_fifo
  inst__maxi_read_req_fifo
  (
    .CLK(CLK),
    .RST(RESETN_inv_buf),
    ._maxi_read_req_fifo_enq(_maxi_read_req_fifo_enq),
    ._maxi_read_req_fifo_wdata(_maxi_read_req_fifo_wdata),
    ._maxi_read_req_fifo_full(_maxi_read_req_fifo_full),
    ._maxi_read_req_fifo_almost_full(_maxi_read_req_fifo_almost_full),
    ._maxi_read_req_fifo_deq(_maxi_read_req_fifo_deq),
    ._maxi_read_req_fifo_rdata(_maxi_read_req_fifo_rdata),
    ._maxi_read_req_fifo_empty(_maxi_read_req_fifo_empty),
    ._maxi_read_req_fifo_almost_empty(_maxi_read_req_fifo_almost_empty)
  );

  reg [4-1:0] count__maxi_read_req_fifo;
  wire [8-1:0] _maxi_read_op_sel_fifo;
  wire [32-1:0] _maxi_read_local_addr_fifo;
  wire [32-1:0] _maxi_read_local_stride_fifo;
  wire [33-1:0] _maxi_read_local_size_fifo;
  wire [32-1:0] _maxi_read_local_blocksize_fifo;
  wire [8-1:0] unpack_read_req_op_sel_30;
  wire [32-1:0] unpack_read_req_local_addr_31;
  wire [32-1:0] unpack_read_req_local_stride_32;
  wire [33-1:0] unpack_read_req_local_size_33;
  wire [32-1:0] unpack_read_req_local_blocksize_34;
  assign unpack_read_req_op_sel_30 = _maxi_read_req_fifo_rdata[136:129];
  assign unpack_read_req_local_addr_31 = _maxi_read_req_fifo_rdata[128:97];
  assign unpack_read_req_local_stride_32 = _maxi_read_req_fifo_rdata[96:65];
  assign unpack_read_req_local_size_33 = _maxi_read_req_fifo_rdata[64:32];
  assign unpack_read_req_local_blocksize_34 = _maxi_read_req_fifo_rdata[31:0];
  assign _maxi_read_op_sel_fifo = unpack_read_req_op_sel_30;
  assign _maxi_read_local_addr_fifo = unpack_read_req_local_addr_31;
  assign _maxi_read_local_stride_fifo = unpack_read_req_local_stride_32;
  assign _maxi_read_local_size_fifo = unpack_read_req_local_size_33;
  assign _maxi_read_local_blocksize_fifo = unpack_read_req_local_blocksize_34;
  reg [8-1:0] _maxi_read_op_sel_buf;
  reg [32-1:0] _maxi_read_local_addr_buf;
  reg [32-1:0] _maxi_read_local_stride_buf;
  reg [33-1:0] _maxi_read_local_size_buf;
  reg [32-1:0] _maxi_read_local_blocksize_buf;
  reg _maxi_read_req_busy;
  reg _maxi_read_data_busy;
  wire _maxi_read_req_idle;
  wire _maxi_read_data_idle;
  wire _maxi_read_idle;
  assign _maxi_read_req_idle = !_maxi_read_start && !_maxi_read_req_busy;
  assign _maxi_read_data_idle = _maxi_read_req_fifo_empty && !_maxi_read_data_busy;
  assign _maxi_read_idle = _maxi_read_req_idle && _maxi_read_data_idle;
  reg _maxi_write_start;
  reg [8-1:0] _maxi_write_op_sel;
  reg [32-1:0] _maxi_write_global_addr;
  reg [33-1:0] _maxi_write_global_size;
  reg [32-1:0] _maxi_write_local_addr;
  reg [32-1:0] _maxi_write_local_stride;
  reg [33-1:0] _maxi_write_local_size;
  reg [32-1:0] _maxi_write_local_blocksize;
  wire _maxi_write_req_fifo_enq;
  wire [137-1:0] _maxi_write_req_fifo_wdata;
  wire _maxi_write_req_fifo_full;
  wire _maxi_write_req_fifo_almost_full;
  wire _maxi_write_req_fifo_deq;
  wire [137-1:0] _maxi_write_req_fifo_rdata;
  wire _maxi_write_req_fifo_empty;
  wire _maxi_write_req_fifo_almost_empty;

  _maxi_write_req_fifo
  inst__maxi_write_req_fifo
  (
    .CLK(CLK),
    .RST(RESETN_inv_buf),
    ._maxi_write_req_fifo_enq(_maxi_write_req_fifo_enq),
    ._maxi_write_req_fifo_wdata(_maxi_write_req_fifo_wdata),
    ._maxi_write_req_fifo_full(_maxi_write_req_fifo_full),
    ._maxi_write_req_fifo_almost_full(_maxi_write_req_fifo_almost_full),
    ._maxi_write_req_fifo_deq(_maxi_write_req_fifo_deq),
    ._maxi_write_req_fifo_rdata(_maxi_write_req_fifo_rdata),
    ._maxi_write_req_fifo_empty(_maxi_write_req_fifo_empty),
    ._maxi_write_req_fifo_almost_empty(_maxi_write_req_fifo_almost_empty)
  );

  reg [4-1:0] count__maxi_write_req_fifo;
  wire [8-1:0] _maxi_write_op_sel_fifo;
  wire [32-1:0] _maxi_write_local_addr_fifo;
  wire [32-1:0] _maxi_write_local_stride_fifo;
  wire [33-1:0] _maxi_write_size_fifo;
  wire [32-1:0] _maxi_write_local_blocksize_fifo;
  wire [8-1:0] unpack_write_req_op_sel_35;
  wire [32-1:0] unpack_write_req_local_addr_36;
  wire [32-1:0] unpack_write_req_local_stride_37;
  wire [33-1:0] unpack_write_req_size_38;
  wire [32-1:0] unpack_write_req_local_blocksize_39;
  assign unpack_write_req_op_sel_35 = _maxi_write_req_fifo_rdata[136:129];
  assign unpack_write_req_local_addr_36 = _maxi_write_req_fifo_rdata[128:97];
  assign unpack_write_req_local_stride_37 = _maxi_write_req_fifo_rdata[96:65];
  assign unpack_write_req_size_38 = _maxi_write_req_fifo_rdata[64:32];
  assign unpack_write_req_local_blocksize_39 = _maxi_write_req_fifo_rdata[31:0];
  assign _maxi_write_op_sel_fifo = unpack_write_req_op_sel_35;
  assign _maxi_write_local_addr_fifo = unpack_write_req_local_addr_36;
  assign _maxi_write_local_stride_fifo = unpack_write_req_local_stride_37;
  assign _maxi_write_size_fifo = unpack_write_req_size_38;
  assign _maxi_write_local_blocksize_fifo = unpack_write_req_local_blocksize_39;
  reg [8-1:0] _maxi_write_op_sel_buf;
  reg [32-1:0] _maxi_write_local_addr_buf;
  reg [32-1:0] _maxi_write_local_stride_buf;
  reg [33-1:0] _maxi_write_size_buf;
  reg [32-1:0] _maxi_write_local_blocksize_buf;
  reg _maxi_write_req_busy;
  reg _maxi_write_data_busy;
  wire _maxi_write_req_idle;
  wire _maxi_write_data_idle;
  wire _maxi_write_idle;
  assign _maxi_write_req_idle = !_maxi_write_start && !_maxi_write_req_busy;
  assign _maxi_write_data_idle = _maxi_write_req_fifo_empty && !_maxi_write_data_busy;
  assign _maxi_write_idle = _maxi_write_req_idle && _maxi_write_data_idle;
  reg [32-1:0] _maxi_global_base_addr;
  assign saxi_bresp = 0;
  assign saxi_rresp = 0;
  reg signed [32-1:0] _saxi_register_0;
  reg signed [32-1:0] _saxi_register_1;
  reg signed [32-1:0] _saxi_register_2;
  reg signed [32-1:0] _saxi_register_3;
  reg signed [32-1:0] _saxi_register_4;
  reg signed [32-1:0] _saxi_register_5;
  reg signed [32-1:0] _saxi_register_6;
  reg signed [32-1:0] _saxi_register_7;
  reg signed [32-1:0] _saxi_register_8;
  reg signed [32-1:0] _saxi_register_9;
  reg signed [32-1:0] _saxi_register_10;
  reg signed [32-1:0] _saxi_register_11;
  reg signed [32-1:0] _saxi_register_12;
  reg signed [32-1:0] _saxi_register_13;
  reg signed [32-1:0] _saxi_register_14;
  reg signed [32-1:0] _saxi_register_15;
  reg signed [32-1:0] _saxi_register_16;
  reg signed [32-1:0] _saxi_register_17;
  reg signed [32-1:0] _saxi_register_18;
  reg signed [32-1:0] _saxi_register_19;
  reg signed [32-1:0] _saxi_register_20;
  reg signed [32-1:0] _saxi_register_21;
  reg signed [32-1:0] _saxi_register_22;
  reg signed [32-1:0] _saxi_register_23;
  reg signed [32-1:0] _saxi_register_24;
  reg signed [32-1:0] _saxi_register_25;
  reg signed [32-1:0] _saxi_register_26;
  reg signed [32-1:0] _saxi_register_27;
  reg signed [32-1:0] _saxi_register_28;
  reg signed [32-1:0] _saxi_register_29;
  reg signed [32-1:0] _saxi_register_30;
  reg signed [32-1:0] _saxi_register_31;
  reg signed [32-1:0] _saxi_register_32;
  reg signed [32-1:0] _saxi_register_33;
  reg signed [32-1:0] _saxi_register_34;
  reg signed [32-1:0] _saxi_register_35;
  reg signed [32-1:0] _saxi_register_36;
  reg _saxi_flag_0;
  reg _saxi_flag_1;
  reg _saxi_flag_2;
  reg _saxi_flag_3;
  reg _saxi_flag_4;
  reg _saxi_flag_5;
  reg _saxi_flag_6;
  reg _saxi_flag_7;
  reg _saxi_flag_8;
  reg _saxi_flag_9;
  reg _saxi_flag_10;
  reg _saxi_flag_11;
  reg _saxi_flag_12;
  reg _saxi_flag_13;
  reg _saxi_flag_14;
  reg _saxi_flag_15;
  reg _saxi_flag_16;
  reg _saxi_flag_17;
  reg _saxi_flag_18;
  reg _saxi_flag_19;
  reg _saxi_flag_20;
  reg _saxi_flag_21;
  reg _saxi_flag_22;
  reg _saxi_flag_23;
  reg _saxi_flag_24;
  reg _saxi_flag_25;
  reg _saxi_flag_26;
  reg _saxi_flag_27;
  reg _saxi_flag_28;
  reg _saxi_flag_29;
  reg _saxi_flag_30;
  reg _saxi_flag_31;
  reg _saxi_flag_32;
  reg _saxi_flag_33;
  reg _saxi_flag_34;
  reg _saxi_flag_35;
  reg _saxi_flag_36;
  reg signed [32-1:0] _saxi_resetval_0;
  reg signed [32-1:0] _saxi_resetval_1;
  reg signed [32-1:0] _saxi_resetval_2;
  reg signed [32-1:0] _saxi_resetval_3;
  reg signed [32-1:0] _saxi_resetval_4;
  reg signed [32-1:0] _saxi_resetval_5;
  reg signed [32-1:0] _saxi_resetval_6;
  reg signed [32-1:0] _saxi_resetval_7;
  reg signed [32-1:0] _saxi_resetval_8;
  reg signed [32-1:0] _saxi_resetval_9;
  reg signed [32-1:0] _saxi_resetval_10;
  reg signed [32-1:0] _saxi_resetval_11;
  reg signed [32-1:0] _saxi_resetval_12;
  reg signed [32-1:0] _saxi_resetval_13;
  reg signed [32-1:0] _saxi_resetval_14;
  reg signed [32-1:0] _saxi_resetval_15;
  reg signed [32-1:0] _saxi_resetval_16;
  reg signed [32-1:0] _saxi_resetval_17;
  reg signed [32-1:0] _saxi_resetval_18;
  reg signed [32-1:0] _saxi_resetval_19;
  reg signed [32-1:0] _saxi_resetval_20;
  reg signed [32-1:0] _saxi_resetval_21;
  reg signed [32-1:0] _saxi_resetval_22;
  reg signed [32-1:0] _saxi_resetval_23;
  reg signed [32-1:0] _saxi_resetval_24;
  reg signed [32-1:0] _saxi_resetval_25;
  reg signed [32-1:0] _saxi_resetval_26;
  reg signed [32-1:0] _saxi_resetval_27;
  reg signed [32-1:0] _saxi_resetval_28;
  reg signed [32-1:0] _saxi_resetval_29;
  reg signed [32-1:0] _saxi_resetval_30;
  reg signed [32-1:0] _saxi_resetval_31;
  reg signed [32-1:0] _saxi_resetval_32;
  reg signed [32-1:0] _saxi_resetval_33;
  reg signed [32-1:0] _saxi_resetval_34;
  reg signed [32-1:0] _saxi_resetval_35;
  reg signed [32-1:0] _saxi_resetval_36;
  localparam _saxi_maskwidth = 6;
  localparam _saxi_mask = { _saxi_maskwidth{ 1'd1 } };
  localparam _saxi_shift = 2;
  reg [32-1:0] _saxi_register_fsm;
  localparam _saxi_register_fsm_init = 0;
  reg [32-1:0] addr_40;
  reg writevalid_41;
  reg readvalid_42;
  reg prev_awvalid_43;
  reg prev_arvalid_44;
  assign saxi_awready = (_saxi_register_fsm == 0) && (!writevalid_41 && !readvalid_42 && !saxi_bvalid && prev_awvalid_43);
  assign saxi_arready = (_saxi_register_fsm == 0) && (!readvalid_42 && !writevalid_41 && prev_arvalid_44 && !prev_awvalid_43);
  reg [_saxi_maskwidth-1:0] axis_maskaddr_45;
  wire signed [32-1:0] axislite_rdata_46;
  assign axislite_rdata_46 = (axis_maskaddr_45 == 0)? _saxi_register_0 : 
                             (axis_maskaddr_45 == 1)? _saxi_register_1 : 
                             (axis_maskaddr_45 == 2)? _saxi_register_2 : 
                             (axis_maskaddr_45 == 3)? _saxi_register_3 : 
                             (axis_maskaddr_45 == 4)? _saxi_register_4 : 
                             (axis_maskaddr_45 == 5)? _saxi_register_5 : 
                             (axis_maskaddr_45 == 6)? _saxi_register_6 : 
                             (axis_maskaddr_45 == 7)? _saxi_register_7 : 
                             (axis_maskaddr_45 == 8)? _saxi_register_8 : 
                             (axis_maskaddr_45 == 9)? _saxi_register_9 : 
                             (axis_maskaddr_45 == 10)? _saxi_register_10 : 
                             (axis_maskaddr_45 == 11)? _saxi_register_11 : 
                             (axis_maskaddr_45 == 12)? _saxi_register_12 : 
                             (axis_maskaddr_45 == 13)? _saxi_register_13 : 
                             (axis_maskaddr_45 == 14)? _saxi_register_14 : 
                             (axis_maskaddr_45 == 15)? _saxi_register_15 : 
                             (axis_maskaddr_45 == 16)? _saxi_register_16 : 
                             (axis_maskaddr_45 == 17)? _saxi_register_17 : 
                             (axis_maskaddr_45 == 18)? _saxi_register_18 : 
                             (axis_maskaddr_45 == 19)? _saxi_register_19 : 
                             (axis_maskaddr_45 == 20)? _saxi_register_20 : 
                             (axis_maskaddr_45 == 21)? _saxi_register_21 : 
                             (axis_maskaddr_45 == 22)? _saxi_register_22 : 
                             (axis_maskaddr_45 == 23)? _saxi_register_23 : 
                             (axis_maskaddr_45 == 24)? _saxi_register_24 : 
                             (axis_maskaddr_45 == 25)? _saxi_register_25 : 
                             (axis_maskaddr_45 == 26)? _saxi_register_26 : 
                             (axis_maskaddr_45 == 27)? _saxi_register_27 : 
                             (axis_maskaddr_45 == 28)? _saxi_register_28 : 
                             (axis_maskaddr_45 == 29)? _saxi_register_29 : 
                             (axis_maskaddr_45 == 30)? _saxi_register_30 : 
                             (axis_maskaddr_45 == 31)? _saxi_register_31 : 
                             (axis_maskaddr_45 == 32)? _saxi_register_32 : 
                             (axis_maskaddr_45 == 33)? _saxi_register_33 : 
                             (axis_maskaddr_45 == 34)? _saxi_register_34 : 
                             (axis_maskaddr_45 == 35)? _saxi_register_35 : 
                             (axis_maskaddr_45 == 36)? _saxi_register_36 : 'hx;
  wire axislite_flag_47;
  assign axislite_flag_47 = (axis_maskaddr_45 == 0)? _saxi_flag_0 : 
                            (axis_maskaddr_45 == 1)? _saxi_flag_1 : 
                            (axis_maskaddr_45 == 2)? _saxi_flag_2 : 
                            (axis_maskaddr_45 == 3)? _saxi_flag_3 : 
                            (axis_maskaddr_45 == 4)? _saxi_flag_4 : 
                            (axis_maskaddr_45 == 5)? _saxi_flag_5 : 
                            (axis_maskaddr_45 == 6)? _saxi_flag_6 : 
                            (axis_maskaddr_45 == 7)? _saxi_flag_7 : 
                            (axis_maskaddr_45 == 8)? _saxi_flag_8 : 
                            (axis_maskaddr_45 == 9)? _saxi_flag_9 : 
                            (axis_maskaddr_45 == 10)? _saxi_flag_10 : 
                            (axis_maskaddr_45 == 11)? _saxi_flag_11 : 
                            (axis_maskaddr_45 == 12)? _saxi_flag_12 : 
                            (axis_maskaddr_45 == 13)? _saxi_flag_13 : 
                            (axis_maskaddr_45 == 14)? _saxi_flag_14 : 
                            (axis_maskaddr_45 == 15)? _saxi_flag_15 : 
                            (axis_maskaddr_45 == 16)? _saxi_flag_16 : 
                            (axis_maskaddr_45 == 17)? _saxi_flag_17 : 
                            (axis_maskaddr_45 == 18)? _saxi_flag_18 : 
                            (axis_maskaddr_45 == 19)? _saxi_flag_19 : 
                            (axis_maskaddr_45 == 20)? _saxi_flag_20 : 
                            (axis_maskaddr_45 == 21)? _saxi_flag_21 : 
                            (axis_maskaddr_45 == 22)? _saxi_flag_22 : 
                            (axis_maskaddr_45 == 23)? _saxi_flag_23 : 
                            (axis_maskaddr_45 == 24)? _saxi_flag_24 : 
                            (axis_maskaddr_45 == 25)? _saxi_flag_25 : 
                            (axis_maskaddr_45 == 26)? _saxi_flag_26 : 
                            (axis_maskaddr_45 == 27)? _saxi_flag_27 : 
                            (axis_maskaddr_45 == 28)? _saxi_flag_28 : 
                            (axis_maskaddr_45 == 29)? _saxi_flag_29 : 
                            (axis_maskaddr_45 == 30)? _saxi_flag_30 : 
                            (axis_maskaddr_45 == 31)? _saxi_flag_31 : 
                            (axis_maskaddr_45 == 32)? _saxi_flag_32 : 
                            (axis_maskaddr_45 == 33)? _saxi_flag_33 : 
                            (axis_maskaddr_45 == 34)? _saxi_flag_34 : 
                            (axis_maskaddr_45 == 35)? _saxi_flag_35 : 
                            (axis_maskaddr_45 == 36)? _saxi_flag_36 : 'hx;
  wire signed [32-1:0] axislite_resetval_48;
  assign axislite_resetval_48 = (axis_maskaddr_45 == 0)? _saxi_resetval_0 : 
                                (axis_maskaddr_45 == 1)? _saxi_resetval_1 : 
                                (axis_maskaddr_45 == 2)? _saxi_resetval_2 : 
                                (axis_maskaddr_45 == 3)? _saxi_resetval_3 : 
                                (axis_maskaddr_45 == 4)? _saxi_resetval_4 : 
                                (axis_maskaddr_45 == 5)? _saxi_resetval_5 : 
                                (axis_maskaddr_45 == 6)? _saxi_resetval_6 : 
                                (axis_maskaddr_45 == 7)? _saxi_resetval_7 : 
                                (axis_maskaddr_45 == 8)? _saxi_resetval_8 : 
                                (axis_maskaddr_45 == 9)? _saxi_resetval_9 : 
                                (axis_maskaddr_45 == 10)? _saxi_resetval_10 : 
                                (axis_maskaddr_45 == 11)? _saxi_resetval_11 : 
                                (axis_maskaddr_45 == 12)? _saxi_resetval_12 : 
                                (axis_maskaddr_45 == 13)? _saxi_resetval_13 : 
                                (axis_maskaddr_45 == 14)? _saxi_resetval_14 : 
                                (axis_maskaddr_45 == 15)? _saxi_resetval_15 : 
                                (axis_maskaddr_45 == 16)? _saxi_resetval_16 : 
                                (axis_maskaddr_45 == 17)? _saxi_resetval_17 : 
                                (axis_maskaddr_45 == 18)? _saxi_resetval_18 : 
                                (axis_maskaddr_45 == 19)? _saxi_resetval_19 : 
                                (axis_maskaddr_45 == 20)? _saxi_resetval_20 : 
                                (axis_maskaddr_45 == 21)? _saxi_resetval_21 : 
                                (axis_maskaddr_45 == 22)? _saxi_resetval_22 : 
                                (axis_maskaddr_45 == 23)? _saxi_resetval_23 : 
                                (axis_maskaddr_45 == 24)? _saxi_resetval_24 : 
                                (axis_maskaddr_45 == 25)? _saxi_resetval_25 : 
                                (axis_maskaddr_45 == 26)? _saxi_resetval_26 : 
                                (axis_maskaddr_45 == 27)? _saxi_resetval_27 : 
                                (axis_maskaddr_45 == 28)? _saxi_resetval_28 : 
                                (axis_maskaddr_45 == 29)? _saxi_resetval_29 : 
                                (axis_maskaddr_45 == 30)? _saxi_resetval_30 : 
                                (axis_maskaddr_45 == 31)? _saxi_resetval_31 : 
                                (axis_maskaddr_45 == 32)? _saxi_resetval_32 : 
                                (axis_maskaddr_45 == 33)? _saxi_resetval_33 : 
                                (axis_maskaddr_45 == 34)? _saxi_resetval_34 : 
                                (axis_maskaddr_45 == 35)? _saxi_resetval_35 : 
                                (axis_maskaddr_45 == 36)? _saxi_resetval_36 : 'hx;
  reg _saxi_rdata_cond_0_1;
  assign saxi_wready = _saxi_register_fsm == 3;
  wire maxi_idle;
  assign maxi_idle = _maxi_write_idle & _maxi_read_idle;
  wire sw_rst_logic;
  assign sw_rst_logic = maxi_idle & _saxi_register_6;
  wire rst_logic;
  assign rst_logic = RESETN_inv_buf | sw_rst_logic;
  reg RST;
  reg _rst_logic_1;
  reg _rst_logic_2;
  wire signed [32-1:0] irq_49;
  assign irq_49 = _saxi_register_9 & _saxi_register_10;
  wire irq_busy;
  assign irq_busy = _saxi_register_5[0];
  reg irq_busy_edge_50;
  wire irq_busy_edge_51;
  assign irq_busy_edge_51 = irq_busy_edge_50 & !irq_busy;
  wire irq_extern;
  assign irq_extern = |_saxi_register_7;
  reg irq_extern_edge_52;
  wire irq_extern_edge_53;
  assign irq_extern_edge_53 = !irq_extern_edge_52 & irq_extern;
  wire [13-1:0] ram_w16_l16384_id0_0_0_addr;
  wire [16-1:0] ram_w16_l16384_id0_0_0_rdata;
  wire [16-1:0] ram_w16_l16384_id0_0_0_wdata;
  wire ram_w16_l16384_id0_0_0_wenable;
  wire ram_w16_l16384_id0_0_0_enable;
  wire [13-1:0] ram_w16_l16384_id0_0_1_addr;
  wire [16-1:0] ram_w16_l16384_id0_0_1_rdata;
  wire [16-1:0] ram_w16_l16384_id0_0_1_wdata;
  wire ram_w16_l16384_id0_0_1_wenable;
  wire ram_w16_l16384_id0_0_1_enable;
  assign ram_w16_l16384_id0_0_0_wdata = 'hx;
  assign ram_w16_l16384_id0_0_0_wenable = 0;

  ram_w16_l16384_id0_0
  inst_ram_w16_l16384_id0_0
  (
    .CLK(CLK),
    .ram_w16_l16384_id0_0_0_addr(ram_w16_l16384_id0_0_0_addr),
    .ram_w16_l16384_id0_0_0_rdata(ram_w16_l16384_id0_0_0_rdata),
    .ram_w16_l16384_id0_0_0_wdata(ram_w16_l16384_id0_0_0_wdata),
    .ram_w16_l16384_id0_0_0_wenable(ram_w16_l16384_id0_0_0_wenable),
    .ram_w16_l16384_id0_0_0_enable(ram_w16_l16384_id0_0_0_enable),
    .ram_w16_l16384_id0_0_1_addr(ram_w16_l16384_id0_0_1_addr),
    .ram_w16_l16384_id0_0_1_rdata(ram_w16_l16384_id0_0_1_rdata),
    .ram_w16_l16384_id0_0_1_wdata(ram_w16_l16384_id0_0_1_wdata),
    .ram_w16_l16384_id0_0_1_wenable(ram_w16_l16384_id0_0_1_wenable),
    .ram_w16_l16384_id0_0_1_enable(ram_w16_l16384_id0_0_1_enable)
  );

  wire [13-1:0] ram_w16_l16384_id0_1_0_addr;
  wire [16-1:0] ram_w16_l16384_id0_1_0_rdata;
  wire [16-1:0] ram_w16_l16384_id0_1_0_wdata;
  wire ram_w16_l16384_id0_1_0_wenable;
  wire ram_w16_l16384_id0_1_0_enable;
  wire [13-1:0] ram_w16_l16384_id0_1_1_addr;
  wire [16-1:0] ram_w16_l16384_id0_1_1_rdata;
  wire [16-1:0] ram_w16_l16384_id0_1_1_wdata;
  wire ram_w16_l16384_id0_1_1_wenable;
  wire ram_w16_l16384_id0_1_1_enable;
  assign ram_w16_l16384_id0_1_0_wdata = 'hx;
  assign ram_w16_l16384_id0_1_0_wenable = 0;

  ram_w16_l16384_id0_1
  inst_ram_w16_l16384_id0_1
  (
    .CLK(CLK),
    .ram_w16_l16384_id0_1_0_addr(ram_w16_l16384_id0_1_0_addr),
    .ram_w16_l16384_id0_1_0_rdata(ram_w16_l16384_id0_1_0_rdata),
    .ram_w16_l16384_id0_1_0_wdata(ram_w16_l16384_id0_1_0_wdata),
    .ram_w16_l16384_id0_1_0_wenable(ram_w16_l16384_id0_1_0_wenable),
    .ram_w16_l16384_id0_1_0_enable(ram_w16_l16384_id0_1_0_enable),
    .ram_w16_l16384_id0_1_1_addr(ram_w16_l16384_id0_1_1_addr),
    .ram_w16_l16384_id0_1_1_rdata(ram_w16_l16384_id0_1_1_rdata),
    .ram_w16_l16384_id0_1_1_wdata(ram_w16_l16384_id0_1_1_wdata),
    .ram_w16_l16384_id0_1_1_wenable(ram_w16_l16384_id0_1_1_wenable),
    .ram_w16_l16384_id0_1_1_enable(ram_w16_l16384_id0_1_1_enable)
  );

  wire [12-1:0] ram_w32_l4096_id0_0_addr;
  wire [32-1:0] ram_w32_l4096_id0_0_rdata;
  wire [32-1:0] ram_w32_l4096_id0_0_wdata;
  wire ram_w32_l4096_id0_0_wenable;
  wire ram_w32_l4096_id0_0_enable;
  wire [12-1:0] ram_w32_l4096_id0_1_addr;
  wire [32-1:0] ram_w32_l4096_id0_1_rdata;
  wire [32-1:0] ram_w32_l4096_id0_1_wdata;
  wire ram_w32_l4096_id0_1_wenable;
  wire ram_w32_l4096_id0_1_enable;
  assign ram_w32_l4096_id0_0_wdata = 'hx;
  assign ram_w32_l4096_id0_0_wenable = 0;

  ram_w32_l4096_id0
  inst_ram_w32_l4096_id0
  (
    .CLK(CLK),
    .ram_w32_l4096_id0_0_addr(ram_w32_l4096_id0_0_addr),
    .ram_w32_l4096_id0_0_rdata(ram_w32_l4096_id0_0_rdata),
    .ram_w32_l4096_id0_0_wdata(ram_w32_l4096_id0_0_wdata),
    .ram_w32_l4096_id0_0_wenable(ram_w32_l4096_id0_0_wenable),
    .ram_w32_l4096_id0_0_enable(ram_w32_l4096_id0_0_enable),
    .ram_w32_l4096_id0_1_addr(ram_w32_l4096_id0_1_addr),
    .ram_w32_l4096_id0_1_rdata(ram_w32_l4096_id0_1_rdata),
    .ram_w32_l4096_id0_1_wdata(ram_w32_l4096_id0_1_wdata),
    .ram_w32_l4096_id0_1_wenable(ram_w32_l4096_id0_1_wenable),
    .ram_w32_l4096_id0_1_enable(ram_w32_l4096_id0_1_enable)
  );

  wire [11-1:0] ram_w16_l4096_id0_0_0_addr;
  wire [16-1:0] ram_w16_l4096_id0_0_0_rdata;
  wire [16-1:0] ram_w16_l4096_id0_0_0_wdata;
  wire ram_w16_l4096_id0_0_0_wenable;
  wire ram_w16_l4096_id0_0_0_enable;
  wire [11-1:0] ram_w16_l4096_id0_0_1_addr;
  wire [16-1:0] ram_w16_l4096_id0_0_1_rdata;
  wire [16-1:0] ram_w16_l4096_id0_0_1_wdata;
  wire ram_w16_l4096_id0_0_1_wenable;
  wire ram_w16_l4096_id0_0_1_enable;
  assign ram_w16_l4096_id0_0_0_wdata = 'hx;
  assign ram_w16_l4096_id0_0_0_wenable = 0;

  ram_w16_l4096_id0_0
  inst_ram_w16_l4096_id0_0
  (
    .CLK(CLK),
    .ram_w16_l4096_id0_0_0_addr(ram_w16_l4096_id0_0_0_addr),
    .ram_w16_l4096_id0_0_0_rdata(ram_w16_l4096_id0_0_0_rdata),
    .ram_w16_l4096_id0_0_0_wdata(ram_w16_l4096_id0_0_0_wdata),
    .ram_w16_l4096_id0_0_0_wenable(ram_w16_l4096_id0_0_0_wenable),
    .ram_w16_l4096_id0_0_0_enable(ram_w16_l4096_id0_0_0_enable),
    .ram_w16_l4096_id0_0_1_addr(ram_w16_l4096_id0_0_1_addr),
    .ram_w16_l4096_id0_0_1_rdata(ram_w16_l4096_id0_0_1_rdata),
    .ram_w16_l4096_id0_0_1_wdata(ram_w16_l4096_id0_0_1_wdata),
    .ram_w16_l4096_id0_0_1_wenable(ram_w16_l4096_id0_0_1_wenable),
    .ram_w16_l4096_id0_0_1_enable(ram_w16_l4096_id0_0_1_enable)
  );

  wire [11-1:0] ram_w16_l4096_id0_1_0_addr;
  wire [16-1:0] ram_w16_l4096_id0_1_0_rdata;
  wire [16-1:0] ram_w16_l4096_id0_1_0_wdata;
  wire ram_w16_l4096_id0_1_0_wenable;
  wire ram_w16_l4096_id0_1_0_enable;
  wire [11-1:0] ram_w16_l4096_id0_1_1_addr;
  wire [16-1:0] ram_w16_l4096_id0_1_1_rdata;
  wire [16-1:0] ram_w16_l4096_id0_1_1_wdata;
  wire ram_w16_l4096_id0_1_1_wenable;
  wire ram_w16_l4096_id0_1_1_enable;
  assign ram_w16_l4096_id0_1_0_wdata = 'hx;
  assign ram_w16_l4096_id0_1_0_wenable = 0;

  ram_w16_l4096_id0_1
  inst_ram_w16_l4096_id0_1
  (
    .CLK(CLK),
    .ram_w16_l4096_id0_1_0_addr(ram_w16_l4096_id0_1_0_addr),
    .ram_w16_l4096_id0_1_0_rdata(ram_w16_l4096_id0_1_0_rdata),
    .ram_w16_l4096_id0_1_0_wdata(ram_w16_l4096_id0_1_0_wdata),
    .ram_w16_l4096_id0_1_0_wenable(ram_w16_l4096_id0_1_0_wenable),
    .ram_w16_l4096_id0_1_0_enable(ram_w16_l4096_id0_1_0_enable),
    .ram_w16_l4096_id0_1_1_addr(ram_w16_l4096_id0_1_1_addr),
    .ram_w16_l4096_id0_1_1_rdata(ram_w16_l4096_id0_1_1_rdata),
    .ram_w16_l4096_id0_1_1_wdata(ram_w16_l4096_id0_1_1_wdata),
    .ram_w16_l4096_id0_1_1_wenable(ram_w16_l4096_id0_1_1_wenable),
    .ram_w16_l4096_id0_1_1_enable(ram_w16_l4096_id0_1_1_enable)
  );

  wire [10-1:0] ram_w32_l1024_id0_0_addr;
  wire [32-1:0] ram_w32_l1024_id0_0_rdata;
  wire [32-1:0] ram_w32_l1024_id0_0_wdata;
  wire ram_w32_l1024_id0_0_wenable;
  wire ram_w32_l1024_id0_0_enable;
  wire [10-1:0] ram_w32_l1024_id0_1_addr;
  wire [32-1:0] ram_w32_l1024_id0_1_rdata;
  wire [32-1:0] ram_w32_l1024_id0_1_wdata;
  wire ram_w32_l1024_id0_1_wenable;
  wire ram_w32_l1024_id0_1_enable;

  ram_w32_l1024_id0
  inst_ram_w32_l1024_id0
  (
    .CLK(CLK),
    .ram_w32_l1024_id0_0_addr(ram_w32_l1024_id0_0_addr),
    .ram_w32_l1024_id0_0_rdata(ram_w32_l1024_id0_0_rdata),
    .ram_w32_l1024_id0_0_wdata(ram_w32_l1024_id0_0_wdata),
    .ram_w32_l1024_id0_0_wenable(ram_w32_l1024_id0_0_wenable),
    .ram_w32_l1024_id0_0_enable(ram_w32_l1024_id0_0_enable),
    .ram_w32_l1024_id0_1_addr(ram_w32_l1024_id0_1_addr),
    .ram_w32_l1024_id0_1_rdata(ram_w32_l1024_id0_1_rdata),
    .ram_w32_l1024_id0_1_wdata(ram_w32_l1024_id0_1_wdata),
    .ram_w32_l1024_id0_1_wenable(ram_w32_l1024_id0_1_wenable),
    .ram_w32_l1024_id0_1_enable(ram_w32_l1024_id0_1_enable)
  );

  wire [9-1:0] ram_w32_l512_id0_0_addr;
  wire [32-1:0] ram_w32_l512_id0_0_rdata;
  wire [32-1:0] ram_w32_l512_id0_0_wdata;
  wire ram_w32_l512_id0_0_wenable;
  wire ram_w32_l512_id0_0_enable;
  wire [9-1:0] ram_w32_l512_id0_1_addr;
  wire [32-1:0] ram_w32_l512_id0_1_rdata;
  wire [32-1:0] ram_w32_l512_id0_1_wdata;
  wire ram_w32_l512_id0_1_wenable;
  wire ram_w32_l512_id0_1_enable;
  assign ram_w32_l512_id0_0_wdata = 'hx;
  assign ram_w32_l512_id0_0_wenable = 0;

  ram_w32_l512_id0
  inst_ram_w32_l512_id0
  (
    .CLK(CLK),
    .ram_w32_l512_id0_0_addr(ram_w32_l512_id0_0_addr),
    .ram_w32_l512_id0_0_rdata(ram_w32_l512_id0_0_rdata),
    .ram_w32_l512_id0_0_wdata(ram_w32_l512_id0_0_wdata),
    .ram_w32_l512_id0_0_wenable(ram_w32_l512_id0_0_wenable),
    .ram_w32_l512_id0_0_enable(ram_w32_l512_id0_0_enable),
    .ram_w32_l512_id0_1_addr(ram_w32_l512_id0_1_addr),
    .ram_w32_l512_id0_1_rdata(ram_w32_l512_id0_1_rdata),
    .ram_w32_l512_id0_1_wdata(ram_w32_l512_id0_1_wdata),
    .ram_w32_l512_id0_1_wenable(ram_w32_l512_id0_1_wenable),
    .ram_w32_l512_id0_1_enable(ram_w32_l512_id0_1_enable)
  );

  wire [9-1:0] ram_w32_l512_id1_0_addr;
  wire [32-1:0] ram_w32_l512_id1_0_rdata;
  wire [32-1:0] ram_w32_l512_id1_0_wdata;
  wire ram_w32_l512_id1_0_wenable;
  wire ram_w32_l512_id1_0_enable;
  wire [9-1:0] ram_w32_l512_id1_1_addr;
  wire [32-1:0] ram_w32_l512_id1_1_rdata;
  wire [32-1:0] ram_w32_l512_id1_1_wdata;
  wire ram_w32_l512_id1_1_wenable;
  wire ram_w32_l512_id1_1_enable;
  assign ram_w32_l512_id1_0_wdata = 'hx;
  assign ram_w32_l512_id1_0_wenable = 0;

  ram_w32_l512_id1
  inst_ram_w32_l512_id1
  (
    .CLK(CLK),
    .ram_w32_l512_id1_0_addr(ram_w32_l512_id1_0_addr),
    .ram_w32_l512_id1_0_rdata(ram_w32_l512_id1_0_rdata),
    .ram_w32_l512_id1_0_wdata(ram_w32_l512_id1_0_wdata),
    .ram_w32_l512_id1_0_wenable(ram_w32_l512_id1_0_wenable),
    .ram_w32_l512_id1_0_enable(ram_w32_l512_id1_0_enable),
    .ram_w32_l512_id1_1_addr(ram_w32_l512_id1_1_addr),
    .ram_w32_l512_id1_1_rdata(ram_w32_l512_id1_1_rdata),
    .ram_w32_l512_id1_1_wdata(ram_w32_l512_id1_1_wdata),
    .ram_w32_l512_id1_1_wenable(ram_w32_l512_id1_1_wenable),
    .ram_w32_l512_id1_1_enable(ram_w32_l512_id1_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id0_0_0_addr;
  wire [16-1:0] ram_w16_l1024_id0_0_0_rdata;
  wire [16-1:0] ram_w16_l1024_id0_0_0_wdata;
  wire ram_w16_l1024_id0_0_0_wenable;
  wire ram_w16_l1024_id0_0_0_enable;
  wire [9-1:0] ram_w16_l1024_id0_0_1_addr;
  wire [16-1:0] ram_w16_l1024_id0_0_1_rdata;
  wire [16-1:0] ram_w16_l1024_id0_0_1_wdata;
  wire ram_w16_l1024_id0_0_1_wenable;
  wire ram_w16_l1024_id0_0_1_enable;
  assign ram_w16_l1024_id0_0_0_wdata = 'hx;
  assign ram_w16_l1024_id0_0_0_wenable = 0;

  ram_w16_l1024_id0_0
  inst_ram_w16_l1024_id0_0
  (
    .CLK(CLK),
    .ram_w16_l1024_id0_0_0_addr(ram_w16_l1024_id0_0_0_addr),
    .ram_w16_l1024_id0_0_0_rdata(ram_w16_l1024_id0_0_0_rdata),
    .ram_w16_l1024_id0_0_0_wdata(ram_w16_l1024_id0_0_0_wdata),
    .ram_w16_l1024_id0_0_0_wenable(ram_w16_l1024_id0_0_0_wenable),
    .ram_w16_l1024_id0_0_0_enable(ram_w16_l1024_id0_0_0_enable),
    .ram_w16_l1024_id0_0_1_addr(ram_w16_l1024_id0_0_1_addr),
    .ram_w16_l1024_id0_0_1_rdata(ram_w16_l1024_id0_0_1_rdata),
    .ram_w16_l1024_id0_0_1_wdata(ram_w16_l1024_id0_0_1_wdata),
    .ram_w16_l1024_id0_0_1_wenable(ram_w16_l1024_id0_0_1_wenable),
    .ram_w16_l1024_id0_0_1_enable(ram_w16_l1024_id0_0_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id0_1_0_addr;
  wire [16-1:0] ram_w16_l1024_id0_1_0_rdata;
  wire [16-1:0] ram_w16_l1024_id0_1_0_wdata;
  wire ram_w16_l1024_id0_1_0_wenable;
  wire ram_w16_l1024_id0_1_0_enable;
  wire [9-1:0] ram_w16_l1024_id0_1_1_addr;
  wire [16-1:0] ram_w16_l1024_id0_1_1_rdata;
  wire [16-1:0] ram_w16_l1024_id0_1_1_wdata;
  wire ram_w16_l1024_id0_1_1_wenable;
  wire ram_w16_l1024_id0_1_1_enable;
  assign ram_w16_l1024_id0_1_0_wdata = 'hx;
  assign ram_w16_l1024_id0_1_0_wenable = 0;

  ram_w16_l1024_id0_1
  inst_ram_w16_l1024_id0_1
  (
    .CLK(CLK),
    .ram_w16_l1024_id0_1_0_addr(ram_w16_l1024_id0_1_0_addr),
    .ram_w16_l1024_id0_1_0_rdata(ram_w16_l1024_id0_1_0_rdata),
    .ram_w16_l1024_id0_1_0_wdata(ram_w16_l1024_id0_1_0_wdata),
    .ram_w16_l1024_id0_1_0_wenable(ram_w16_l1024_id0_1_0_wenable),
    .ram_w16_l1024_id0_1_0_enable(ram_w16_l1024_id0_1_0_enable),
    .ram_w16_l1024_id0_1_1_addr(ram_w16_l1024_id0_1_1_addr),
    .ram_w16_l1024_id0_1_1_rdata(ram_w16_l1024_id0_1_1_rdata),
    .ram_w16_l1024_id0_1_1_wdata(ram_w16_l1024_id0_1_1_wdata),
    .ram_w16_l1024_id0_1_1_wenable(ram_w16_l1024_id0_1_1_wenable),
    .ram_w16_l1024_id0_1_1_enable(ram_w16_l1024_id0_1_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id1_0_0_addr;
  wire [16-1:0] ram_w16_l1024_id1_0_0_rdata;
  wire [16-1:0] ram_w16_l1024_id1_0_0_wdata;
  wire ram_w16_l1024_id1_0_0_wenable;
  wire ram_w16_l1024_id1_0_0_enable;
  wire [9-1:0] ram_w16_l1024_id1_0_1_addr;
  wire [16-1:0] ram_w16_l1024_id1_0_1_rdata;
  wire [16-1:0] ram_w16_l1024_id1_0_1_wdata;
  wire ram_w16_l1024_id1_0_1_wenable;
  wire ram_w16_l1024_id1_0_1_enable;
  assign ram_w16_l1024_id1_0_0_wdata = 'hx;
  assign ram_w16_l1024_id1_0_0_wenable = 0;

  ram_w16_l1024_id1_0
  inst_ram_w16_l1024_id1_0
  (
    .CLK(CLK),
    .ram_w16_l1024_id1_0_0_addr(ram_w16_l1024_id1_0_0_addr),
    .ram_w16_l1024_id1_0_0_rdata(ram_w16_l1024_id1_0_0_rdata),
    .ram_w16_l1024_id1_0_0_wdata(ram_w16_l1024_id1_0_0_wdata),
    .ram_w16_l1024_id1_0_0_wenable(ram_w16_l1024_id1_0_0_wenable),
    .ram_w16_l1024_id1_0_0_enable(ram_w16_l1024_id1_0_0_enable),
    .ram_w16_l1024_id1_0_1_addr(ram_w16_l1024_id1_0_1_addr),
    .ram_w16_l1024_id1_0_1_rdata(ram_w16_l1024_id1_0_1_rdata),
    .ram_w16_l1024_id1_0_1_wdata(ram_w16_l1024_id1_0_1_wdata),
    .ram_w16_l1024_id1_0_1_wenable(ram_w16_l1024_id1_0_1_wenable),
    .ram_w16_l1024_id1_0_1_enable(ram_w16_l1024_id1_0_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id1_1_0_addr;
  wire [16-1:0] ram_w16_l1024_id1_1_0_rdata;
  wire [16-1:0] ram_w16_l1024_id1_1_0_wdata;
  wire ram_w16_l1024_id1_1_0_wenable;
  wire ram_w16_l1024_id1_1_0_enable;
  wire [9-1:0] ram_w16_l1024_id1_1_1_addr;
  wire [16-1:0] ram_w16_l1024_id1_1_1_rdata;
  wire [16-1:0] ram_w16_l1024_id1_1_1_wdata;
  wire ram_w16_l1024_id1_1_1_wenable;
  wire ram_w16_l1024_id1_1_1_enable;
  assign ram_w16_l1024_id1_1_0_wdata = 'hx;
  assign ram_w16_l1024_id1_1_0_wenable = 0;

  ram_w16_l1024_id1_1
  inst_ram_w16_l1024_id1_1
  (
    .CLK(CLK),
    .ram_w16_l1024_id1_1_0_addr(ram_w16_l1024_id1_1_0_addr),
    .ram_w16_l1024_id1_1_0_rdata(ram_w16_l1024_id1_1_0_rdata),
    .ram_w16_l1024_id1_1_0_wdata(ram_w16_l1024_id1_1_0_wdata),
    .ram_w16_l1024_id1_1_0_wenable(ram_w16_l1024_id1_1_0_wenable),
    .ram_w16_l1024_id1_1_0_enable(ram_w16_l1024_id1_1_0_enable),
    .ram_w16_l1024_id1_1_1_addr(ram_w16_l1024_id1_1_1_addr),
    .ram_w16_l1024_id1_1_1_rdata(ram_w16_l1024_id1_1_1_rdata),
    .ram_w16_l1024_id1_1_1_wdata(ram_w16_l1024_id1_1_1_wdata),
    .ram_w16_l1024_id1_1_1_wenable(ram_w16_l1024_id1_1_1_wenable),
    .ram_w16_l1024_id1_1_1_enable(ram_w16_l1024_id1_1_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id2_0_0_addr;
  wire [16-1:0] ram_w16_l1024_id2_0_0_rdata;
  wire [16-1:0] ram_w16_l1024_id2_0_0_wdata;
  wire ram_w16_l1024_id2_0_0_wenable;
  wire ram_w16_l1024_id2_0_0_enable;
  wire [9-1:0] ram_w16_l1024_id2_0_1_addr;
  wire [16-1:0] ram_w16_l1024_id2_0_1_rdata;
  wire [16-1:0] ram_w16_l1024_id2_0_1_wdata;
  wire ram_w16_l1024_id2_0_1_wenable;
  wire ram_w16_l1024_id2_0_1_enable;
  assign ram_w16_l1024_id2_0_0_wdata = 'hx;
  assign ram_w16_l1024_id2_0_0_wenable = 0;

  ram_w16_l1024_id2_0
  inst_ram_w16_l1024_id2_0
  (
    .CLK(CLK),
    .ram_w16_l1024_id2_0_0_addr(ram_w16_l1024_id2_0_0_addr),
    .ram_w16_l1024_id2_0_0_rdata(ram_w16_l1024_id2_0_0_rdata),
    .ram_w16_l1024_id2_0_0_wdata(ram_w16_l1024_id2_0_0_wdata),
    .ram_w16_l1024_id2_0_0_wenable(ram_w16_l1024_id2_0_0_wenable),
    .ram_w16_l1024_id2_0_0_enable(ram_w16_l1024_id2_0_0_enable),
    .ram_w16_l1024_id2_0_1_addr(ram_w16_l1024_id2_0_1_addr),
    .ram_w16_l1024_id2_0_1_rdata(ram_w16_l1024_id2_0_1_rdata),
    .ram_w16_l1024_id2_0_1_wdata(ram_w16_l1024_id2_0_1_wdata),
    .ram_w16_l1024_id2_0_1_wenable(ram_w16_l1024_id2_0_1_wenable),
    .ram_w16_l1024_id2_0_1_enable(ram_w16_l1024_id2_0_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id2_1_0_addr;
  wire [16-1:0] ram_w16_l1024_id2_1_0_rdata;
  wire [16-1:0] ram_w16_l1024_id2_1_0_wdata;
  wire ram_w16_l1024_id2_1_0_wenable;
  wire ram_w16_l1024_id2_1_0_enable;
  wire [9-1:0] ram_w16_l1024_id2_1_1_addr;
  wire [16-1:0] ram_w16_l1024_id2_1_1_rdata;
  wire [16-1:0] ram_w16_l1024_id2_1_1_wdata;
  wire ram_w16_l1024_id2_1_1_wenable;
  wire ram_w16_l1024_id2_1_1_enable;
  assign ram_w16_l1024_id2_1_0_wdata = 'hx;
  assign ram_w16_l1024_id2_1_0_wenable = 0;

  ram_w16_l1024_id2_1
  inst_ram_w16_l1024_id2_1
  (
    .CLK(CLK),
    .ram_w16_l1024_id2_1_0_addr(ram_w16_l1024_id2_1_0_addr),
    .ram_w16_l1024_id2_1_0_rdata(ram_w16_l1024_id2_1_0_rdata),
    .ram_w16_l1024_id2_1_0_wdata(ram_w16_l1024_id2_1_0_wdata),
    .ram_w16_l1024_id2_1_0_wenable(ram_w16_l1024_id2_1_0_wenable),
    .ram_w16_l1024_id2_1_0_enable(ram_w16_l1024_id2_1_0_enable),
    .ram_w16_l1024_id2_1_1_addr(ram_w16_l1024_id2_1_1_addr),
    .ram_w16_l1024_id2_1_1_rdata(ram_w16_l1024_id2_1_1_rdata),
    .ram_w16_l1024_id2_1_1_wdata(ram_w16_l1024_id2_1_1_wdata),
    .ram_w16_l1024_id2_1_1_wenable(ram_w16_l1024_id2_1_1_wenable),
    .ram_w16_l1024_id2_1_1_enable(ram_w16_l1024_id2_1_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id3_0_0_addr;
  wire [16-1:0] ram_w16_l1024_id3_0_0_rdata;
  wire [16-1:0] ram_w16_l1024_id3_0_0_wdata;
  wire ram_w16_l1024_id3_0_0_wenable;
  wire ram_w16_l1024_id3_0_0_enable;
  wire [9-1:0] ram_w16_l1024_id3_0_1_addr;
  wire [16-1:0] ram_w16_l1024_id3_0_1_rdata;
  wire [16-1:0] ram_w16_l1024_id3_0_1_wdata;
  wire ram_w16_l1024_id3_0_1_wenable;
  wire ram_w16_l1024_id3_0_1_enable;
  assign ram_w16_l1024_id3_0_0_wdata = 'hx;
  assign ram_w16_l1024_id3_0_0_wenable = 0;

  ram_w16_l1024_id3_0
  inst_ram_w16_l1024_id3_0
  (
    .CLK(CLK),
    .ram_w16_l1024_id3_0_0_addr(ram_w16_l1024_id3_0_0_addr),
    .ram_w16_l1024_id3_0_0_rdata(ram_w16_l1024_id3_0_0_rdata),
    .ram_w16_l1024_id3_0_0_wdata(ram_w16_l1024_id3_0_0_wdata),
    .ram_w16_l1024_id3_0_0_wenable(ram_w16_l1024_id3_0_0_wenable),
    .ram_w16_l1024_id3_0_0_enable(ram_w16_l1024_id3_0_0_enable),
    .ram_w16_l1024_id3_0_1_addr(ram_w16_l1024_id3_0_1_addr),
    .ram_w16_l1024_id3_0_1_rdata(ram_w16_l1024_id3_0_1_rdata),
    .ram_w16_l1024_id3_0_1_wdata(ram_w16_l1024_id3_0_1_wdata),
    .ram_w16_l1024_id3_0_1_wenable(ram_w16_l1024_id3_0_1_wenable),
    .ram_w16_l1024_id3_0_1_enable(ram_w16_l1024_id3_0_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id3_1_0_addr;
  wire [16-1:0] ram_w16_l1024_id3_1_0_rdata;
  wire [16-1:0] ram_w16_l1024_id3_1_0_wdata;
  wire ram_w16_l1024_id3_1_0_wenable;
  wire ram_w16_l1024_id3_1_0_enable;
  wire [9-1:0] ram_w16_l1024_id3_1_1_addr;
  wire [16-1:0] ram_w16_l1024_id3_1_1_rdata;
  wire [16-1:0] ram_w16_l1024_id3_1_1_wdata;
  wire ram_w16_l1024_id3_1_1_wenable;
  wire ram_w16_l1024_id3_1_1_enable;
  assign ram_w16_l1024_id3_1_0_wdata = 'hx;
  assign ram_w16_l1024_id3_1_0_wenable = 0;

  ram_w16_l1024_id3_1
  inst_ram_w16_l1024_id3_1
  (
    .CLK(CLK),
    .ram_w16_l1024_id3_1_0_addr(ram_w16_l1024_id3_1_0_addr),
    .ram_w16_l1024_id3_1_0_rdata(ram_w16_l1024_id3_1_0_rdata),
    .ram_w16_l1024_id3_1_0_wdata(ram_w16_l1024_id3_1_0_wdata),
    .ram_w16_l1024_id3_1_0_wenable(ram_w16_l1024_id3_1_0_wenable),
    .ram_w16_l1024_id3_1_0_enable(ram_w16_l1024_id3_1_0_enable),
    .ram_w16_l1024_id3_1_1_addr(ram_w16_l1024_id3_1_1_addr),
    .ram_w16_l1024_id3_1_1_rdata(ram_w16_l1024_id3_1_1_rdata),
    .ram_w16_l1024_id3_1_1_wdata(ram_w16_l1024_id3_1_1_wdata),
    .ram_w16_l1024_id3_1_1_wenable(ram_w16_l1024_id3_1_1_wenable),
    .ram_w16_l1024_id3_1_1_enable(ram_w16_l1024_id3_1_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id4_0_0_addr;
  wire [16-1:0] ram_w16_l1024_id4_0_0_rdata;
  wire [16-1:0] ram_w16_l1024_id4_0_0_wdata;
  wire ram_w16_l1024_id4_0_0_wenable;
  wire ram_w16_l1024_id4_0_0_enable;
  wire [9-1:0] ram_w16_l1024_id4_0_1_addr;
  wire [16-1:0] ram_w16_l1024_id4_0_1_rdata;
  wire [16-1:0] ram_w16_l1024_id4_0_1_wdata;
  wire ram_w16_l1024_id4_0_1_wenable;
  wire ram_w16_l1024_id4_0_1_enable;
  assign ram_w16_l1024_id4_0_0_wdata = 'hx;
  assign ram_w16_l1024_id4_0_0_wenable = 0;

  ram_w16_l1024_id4_0
  inst_ram_w16_l1024_id4_0
  (
    .CLK(CLK),
    .ram_w16_l1024_id4_0_0_addr(ram_w16_l1024_id4_0_0_addr),
    .ram_w16_l1024_id4_0_0_rdata(ram_w16_l1024_id4_0_0_rdata),
    .ram_w16_l1024_id4_0_0_wdata(ram_w16_l1024_id4_0_0_wdata),
    .ram_w16_l1024_id4_0_0_wenable(ram_w16_l1024_id4_0_0_wenable),
    .ram_w16_l1024_id4_0_0_enable(ram_w16_l1024_id4_0_0_enable),
    .ram_w16_l1024_id4_0_1_addr(ram_w16_l1024_id4_0_1_addr),
    .ram_w16_l1024_id4_0_1_rdata(ram_w16_l1024_id4_0_1_rdata),
    .ram_w16_l1024_id4_0_1_wdata(ram_w16_l1024_id4_0_1_wdata),
    .ram_w16_l1024_id4_0_1_wenable(ram_w16_l1024_id4_0_1_wenable),
    .ram_w16_l1024_id4_0_1_enable(ram_w16_l1024_id4_0_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id4_1_0_addr;
  wire [16-1:0] ram_w16_l1024_id4_1_0_rdata;
  wire [16-1:0] ram_w16_l1024_id4_1_0_wdata;
  wire ram_w16_l1024_id4_1_0_wenable;
  wire ram_w16_l1024_id4_1_0_enable;
  wire [9-1:0] ram_w16_l1024_id4_1_1_addr;
  wire [16-1:0] ram_w16_l1024_id4_1_1_rdata;
  wire [16-1:0] ram_w16_l1024_id4_1_1_wdata;
  wire ram_w16_l1024_id4_1_1_wenable;
  wire ram_w16_l1024_id4_1_1_enable;
  assign ram_w16_l1024_id4_1_0_wdata = 'hx;
  assign ram_w16_l1024_id4_1_0_wenable = 0;

  ram_w16_l1024_id4_1
  inst_ram_w16_l1024_id4_1
  (
    .CLK(CLK),
    .ram_w16_l1024_id4_1_0_addr(ram_w16_l1024_id4_1_0_addr),
    .ram_w16_l1024_id4_1_0_rdata(ram_w16_l1024_id4_1_0_rdata),
    .ram_w16_l1024_id4_1_0_wdata(ram_w16_l1024_id4_1_0_wdata),
    .ram_w16_l1024_id4_1_0_wenable(ram_w16_l1024_id4_1_0_wenable),
    .ram_w16_l1024_id4_1_0_enable(ram_w16_l1024_id4_1_0_enable),
    .ram_w16_l1024_id4_1_1_addr(ram_w16_l1024_id4_1_1_addr),
    .ram_w16_l1024_id4_1_1_rdata(ram_w16_l1024_id4_1_1_rdata),
    .ram_w16_l1024_id4_1_1_wdata(ram_w16_l1024_id4_1_1_wdata),
    .ram_w16_l1024_id4_1_1_wenable(ram_w16_l1024_id4_1_1_wenable),
    .ram_w16_l1024_id4_1_1_enable(ram_w16_l1024_id4_1_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id5_0_0_addr;
  wire [16-1:0] ram_w16_l1024_id5_0_0_rdata;
  wire [16-1:0] ram_w16_l1024_id5_0_0_wdata;
  wire ram_w16_l1024_id5_0_0_wenable;
  wire ram_w16_l1024_id5_0_0_enable;
  wire [9-1:0] ram_w16_l1024_id5_0_1_addr;
  wire [16-1:0] ram_w16_l1024_id5_0_1_rdata;
  wire [16-1:0] ram_w16_l1024_id5_0_1_wdata;
  wire ram_w16_l1024_id5_0_1_wenable;
  wire ram_w16_l1024_id5_0_1_enable;
  assign ram_w16_l1024_id5_0_0_wdata = 'hx;
  assign ram_w16_l1024_id5_0_0_wenable = 0;

  ram_w16_l1024_id5_0
  inst_ram_w16_l1024_id5_0
  (
    .CLK(CLK),
    .ram_w16_l1024_id5_0_0_addr(ram_w16_l1024_id5_0_0_addr),
    .ram_w16_l1024_id5_0_0_rdata(ram_w16_l1024_id5_0_0_rdata),
    .ram_w16_l1024_id5_0_0_wdata(ram_w16_l1024_id5_0_0_wdata),
    .ram_w16_l1024_id5_0_0_wenable(ram_w16_l1024_id5_0_0_wenable),
    .ram_w16_l1024_id5_0_0_enable(ram_w16_l1024_id5_0_0_enable),
    .ram_w16_l1024_id5_0_1_addr(ram_w16_l1024_id5_0_1_addr),
    .ram_w16_l1024_id5_0_1_rdata(ram_w16_l1024_id5_0_1_rdata),
    .ram_w16_l1024_id5_0_1_wdata(ram_w16_l1024_id5_0_1_wdata),
    .ram_w16_l1024_id5_0_1_wenable(ram_w16_l1024_id5_0_1_wenable),
    .ram_w16_l1024_id5_0_1_enable(ram_w16_l1024_id5_0_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id5_1_0_addr;
  wire [16-1:0] ram_w16_l1024_id5_1_0_rdata;
  wire [16-1:0] ram_w16_l1024_id5_1_0_wdata;
  wire ram_w16_l1024_id5_1_0_wenable;
  wire ram_w16_l1024_id5_1_0_enable;
  wire [9-1:0] ram_w16_l1024_id5_1_1_addr;
  wire [16-1:0] ram_w16_l1024_id5_1_1_rdata;
  wire [16-1:0] ram_w16_l1024_id5_1_1_wdata;
  wire ram_w16_l1024_id5_1_1_wenable;
  wire ram_w16_l1024_id5_1_1_enable;
  assign ram_w16_l1024_id5_1_0_wdata = 'hx;
  assign ram_w16_l1024_id5_1_0_wenable = 0;

  ram_w16_l1024_id5_1
  inst_ram_w16_l1024_id5_1
  (
    .CLK(CLK),
    .ram_w16_l1024_id5_1_0_addr(ram_w16_l1024_id5_1_0_addr),
    .ram_w16_l1024_id5_1_0_rdata(ram_w16_l1024_id5_1_0_rdata),
    .ram_w16_l1024_id5_1_0_wdata(ram_w16_l1024_id5_1_0_wdata),
    .ram_w16_l1024_id5_1_0_wenable(ram_w16_l1024_id5_1_0_wenable),
    .ram_w16_l1024_id5_1_0_enable(ram_w16_l1024_id5_1_0_enable),
    .ram_w16_l1024_id5_1_1_addr(ram_w16_l1024_id5_1_1_addr),
    .ram_w16_l1024_id5_1_1_rdata(ram_w16_l1024_id5_1_1_rdata),
    .ram_w16_l1024_id5_1_1_wdata(ram_w16_l1024_id5_1_1_wdata),
    .ram_w16_l1024_id5_1_1_wenable(ram_w16_l1024_id5_1_1_wenable),
    .ram_w16_l1024_id5_1_1_enable(ram_w16_l1024_id5_1_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id6_0_0_addr;
  wire [16-1:0] ram_w16_l1024_id6_0_0_rdata;
  wire [16-1:0] ram_w16_l1024_id6_0_0_wdata;
  wire ram_w16_l1024_id6_0_0_wenable;
  wire ram_w16_l1024_id6_0_0_enable;
  wire [9-1:0] ram_w16_l1024_id6_0_1_addr;
  wire [16-1:0] ram_w16_l1024_id6_0_1_rdata;
  wire [16-1:0] ram_w16_l1024_id6_0_1_wdata;
  wire ram_w16_l1024_id6_0_1_wenable;
  wire ram_w16_l1024_id6_0_1_enable;
  assign ram_w16_l1024_id6_0_0_wdata = 'hx;
  assign ram_w16_l1024_id6_0_0_wenable = 0;

  ram_w16_l1024_id6_0
  inst_ram_w16_l1024_id6_0
  (
    .CLK(CLK),
    .ram_w16_l1024_id6_0_0_addr(ram_w16_l1024_id6_0_0_addr),
    .ram_w16_l1024_id6_0_0_rdata(ram_w16_l1024_id6_0_0_rdata),
    .ram_w16_l1024_id6_0_0_wdata(ram_w16_l1024_id6_0_0_wdata),
    .ram_w16_l1024_id6_0_0_wenable(ram_w16_l1024_id6_0_0_wenable),
    .ram_w16_l1024_id6_0_0_enable(ram_w16_l1024_id6_0_0_enable),
    .ram_w16_l1024_id6_0_1_addr(ram_w16_l1024_id6_0_1_addr),
    .ram_w16_l1024_id6_0_1_rdata(ram_w16_l1024_id6_0_1_rdata),
    .ram_w16_l1024_id6_0_1_wdata(ram_w16_l1024_id6_0_1_wdata),
    .ram_w16_l1024_id6_0_1_wenable(ram_w16_l1024_id6_0_1_wenable),
    .ram_w16_l1024_id6_0_1_enable(ram_w16_l1024_id6_0_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id6_1_0_addr;
  wire [16-1:0] ram_w16_l1024_id6_1_0_rdata;
  wire [16-1:0] ram_w16_l1024_id6_1_0_wdata;
  wire ram_w16_l1024_id6_1_0_wenable;
  wire ram_w16_l1024_id6_1_0_enable;
  wire [9-1:0] ram_w16_l1024_id6_1_1_addr;
  wire [16-1:0] ram_w16_l1024_id6_1_1_rdata;
  wire [16-1:0] ram_w16_l1024_id6_1_1_wdata;
  wire ram_w16_l1024_id6_1_1_wenable;
  wire ram_w16_l1024_id6_1_1_enable;
  assign ram_w16_l1024_id6_1_0_wdata = 'hx;
  assign ram_w16_l1024_id6_1_0_wenable = 0;

  ram_w16_l1024_id6_1
  inst_ram_w16_l1024_id6_1
  (
    .CLK(CLK),
    .ram_w16_l1024_id6_1_0_addr(ram_w16_l1024_id6_1_0_addr),
    .ram_w16_l1024_id6_1_0_rdata(ram_w16_l1024_id6_1_0_rdata),
    .ram_w16_l1024_id6_1_0_wdata(ram_w16_l1024_id6_1_0_wdata),
    .ram_w16_l1024_id6_1_0_wenable(ram_w16_l1024_id6_1_0_wenable),
    .ram_w16_l1024_id6_1_0_enable(ram_w16_l1024_id6_1_0_enable),
    .ram_w16_l1024_id6_1_1_addr(ram_w16_l1024_id6_1_1_addr),
    .ram_w16_l1024_id6_1_1_rdata(ram_w16_l1024_id6_1_1_rdata),
    .ram_w16_l1024_id6_1_1_wdata(ram_w16_l1024_id6_1_1_wdata),
    .ram_w16_l1024_id6_1_1_wenable(ram_w16_l1024_id6_1_1_wenable),
    .ram_w16_l1024_id6_1_1_enable(ram_w16_l1024_id6_1_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id7_0_0_addr;
  wire [16-1:0] ram_w16_l1024_id7_0_0_rdata;
  wire [16-1:0] ram_w16_l1024_id7_0_0_wdata;
  wire ram_w16_l1024_id7_0_0_wenable;
  wire ram_w16_l1024_id7_0_0_enable;
  wire [9-1:0] ram_w16_l1024_id7_0_1_addr;
  wire [16-1:0] ram_w16_l1024_id7_0_1_rdata;
  wire [16-1:0] ram_w16_l1024_id7_0_1_wdata;
  wire ram_w16_l1024_id7_0_1_wenable;
  wire ram_w16_l1024_id7_0_1_enable;
  assign ram_w16_l1024_id7_0_0_wdata = 'hx;
  assign ram_w16_l1024_id7_0_0_wenable = 0;

  ram_w16_l1024_id7_0
  inst_ram_w16_l1024_id7_0
  (
    .CLK(CLK),
    .ram_w16_l1024_id7_0_0_addr(ram_w16_l1024_id7_0_0_addr),
    .ram_w16_l1024_id7_0_0_rdata(ram_w16_l1024_id7_0_0_rdata),
    .ram_w16_l1024_id7_0_0_wdata(ram_w16_l1024_id7_0_0_wdata),
    .ram_w16_l1024_id7_0_0_wenable(ram_w16_l1024_id7_0_0_wenable),
    .ram_w16_l1024_id7_0_0_enable(ram_w16_l1024_id7_0_0_enable),
    .ram_w16_l1024_id7_0_1_addr(ram_w16_l1024_id7_0_1_addr),
    .ram_w16_l1024_id7_0_1_rdata(ram_w16_l1024_id7_0_1_rdata),
    .ram_w16_l1024_id7_0_1_wdata(ram_w16_l1024_id7_0_1_wdata),
    .ram_w16_l1024_id7_0_1_wenable(ram_w16_l1024_id7_0_1_wenable),
    .ram_w16_l1024_id7_0_1_enable(ram_w16_l1024_id7_0_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id7_1_0_addr;
  wire [16-1:0] ram_w16_l1024_id7_1_0_rdata;
  wire [16-1:0] ram_w16_l1024_id7_1_0_wdata;
  wire ram_w16_l1024_id7_1_0_wenable;
  wire ram_w16_l1024_id7_1_0_enable;
  wire [9-1:0] ram_w16_l1024_id7_1_1_addr;
  wire [16-1:0] ram_w16_l1024_id7_1_1_rdata;
  wire [16-1:0] ram_w16_l1024_id7_1_1_wdata;
  wire ram_w16_l1024_id7_1_1_wenable;
  wire ram_w16_l1024_id7_1_1_enable;
  assign ram_w16_l1024_id7_1_0_wdata = 'hx;
  assign ram_w16_l1024_id7_1_0_wenable = 0;

  ram_w16_l1024_id7_1
  inst_ram_w16_l1024_id7_1
  (
    .CLK(CLK),
    .ram_w16_l1024_id7_1_0_addr(ram_w16_l1024_id7_1_0_addr),
    .ram_w16_l1024_id7_1_0_rdata(ram_w16_l1024_id7_1_0_rdata),
    .ram_w16_l1024_id7_1_0_wdata(ram_w16_l1024_id7_1_0_wdata),
    .ram_w16_l1024_id7_1_0_wenable(ram_w16_l1024_id7_1_0_wenable),
    .ram_w16_l1024_id7_1_0_enable(ram_w16_l1024_id7_1_0_enable),
    .ram_w16_l1024_id7_1_1_addr(ram_w16_l1024_id7_1_1_addr),
    .ram_w16_l1024_id7_1_1_rdata(ram_w16_l1024_id7_1_1_rdata),
    .ram_w16_l1024_id7_1_1_wdata(ram_w16_l1024_id7_1_1_wdata),
    .ram_w16_l1024_id7_1_1_wenable(ram_w16_l1024_id7_1_1_wenable),
    .ram_w16_l1024_id7_1_1_enable(ram_w16_l1024_id7_1_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id8_0_0_addr;
  wire [16-1:0] ram_w16_l1024_id8_0_0_rdata;
  wire [16-1:0] ram_w16_l1024_id8_0_0_wdata;
  wire ram_w16_l1024_id8_0_0_wenable;
  wire ram_w16_l1024_id8_0_0_enable;
  wire [9-1:0] ram_w16_l1024_id8_0_1_addr;
  wire [16-1:0] ram_w16_l1024_id8_0_1_rdata;
  wire [16-1:0] ram_w16_l1024_id8_0_1_wdata;
  wire ram_w16_l1024_id8_0_1_wenable;
  wire ram_w16_l1024_id8_0_1_enable;
  assign ram_w16_l1024_id8_0_0_wdata = 'hx;
  assign ram_w16_l1024_id8_0_0_wenable = 0;

  ram_w16_l1024_id8_0
  inst_ram_w16_l1024_id8_0
  (
    .CLK(CLK),
    .ram_w16_l1024_id8_0_0_addr(ram_w16_l1024_id8_0_0_addr),
    .ram_w16_l1024_id8_0_0_rdata(ram_w16_l1024_id8_0_0_rdata),
    .ram_w16_l1024_id8_0_0_wdata(ram_w16_l1024_id8_0_0_wdata),
    .ram_w16_l1024_id8_0_0_wenable(ram_w16_l1024_id8_0_0_wenable),
    .ram_w16_l1024_id8_0_0_enable(ram_w16_l1024_id8_0_0_enable),
    .ram_w16_l1024_id8_0_1_addr(ram_w16_l1024_id8_0_1_addr),
    .ram_w16_l1024_id8_0_1_rdata(ram_w16_l1024_id8_0_1_rdata),
    .ram_w16_l1024_id8_0_1_wdata(ram_w16_l1024_id8_0_1_wdata),
    .ram_w16_l1024_id8_0_1_wenable(ram_w16_l1024_id8_0_1_wenable),
    .ram_w16_l1024_id8_0_1_enable(ram_w16_l1024_id8_0_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id8_1_0_addr;
  wire [16-1:0] ram_w16_l1024_id8_1_0_rdata;
  wire [16-1:0] ram_w16_l1024_id8_1_0_wdata;
  wire ram_w16_l1024_id8_1_0_wenable;
  wire ram_w16_l1024_id8_1_0_enable;
  wire [9-1:0] ram_w16_l1024_id8_1_1_addr;
  wire [16-1:0] ram_w16_l1024_id8_1_1_rdata;
  wire [16-1:0] ram_w16_l1024_id8_1_1_wdata;
  wire ram_w16_l1024_id8_1_1_wenable;
  wire ram_w16_l1024_id8_1_1_enable;
  assign ram_w16_l1024_id8_1_0_wdata = 'hx;
  assign ram_w16_l1024_id8_1_0_wenable = 0;

  ram_w16_l1024_id8_1
  inst_ram_w16_l1024_id8_1
  (
    .CLK(CLK),
    .ram_w16_l1024_id8_1_0_addr(ram_w16_l1024_id8_1_0_addr),
    .ram_w16_l1024_id8_1_0_rdata(ram_w16_l1024_id8_1_0_rdata),
    .ram_w16_l1024_id8_1_0_wdata(ram_w16_l1024_id8_1_0_wdata),
    .ram_w16_l1024_id8_1_0_wenable(ram_w16_l1024_id8_1_0_wenable),
    .ram_w16_l1024_id8_1_0_enable(ram_w16_l1024_id8_1_0_enable),
    .ram_w16_l1024_id8_1_1_addr(ram_w16_l1024_id8_1_1_addr),
    .ram_w16_l1024_id8_1_1_rdata(ram_w16_l1024_id8_1_1_rdata),
    .ram_w16_l1024_id8_1_1_wdata(ram_w16_l1024_id8_1_1_wdata),
    .ram_w16_l1024_id8_1_1_wenable(ram_w16_l1024_id8_1_1_wenable),
    .ram_w16_l1024_id8_1_1_enable(ram_w16_l1024_id8_1_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id9_0_0_addr;
  wire [16-1:0] ram_w16_l1024_id9_0_0_rdata;
  wire [16-1:0] ram_w16_l1024_id9_0_0_wdata;
  wire ram_w16_l1024_id9_0_0_wenable;
  wire ram_w16_l1024_id9_0_0_enable;
  wire [9-1:0] ram_w16_l1024_id9_0_1_addr;
  wire [16-1:0] ram_w16_l1024_id9_0_1_rdata;
  wire [16-1:0] ram_w16_l1024_id9_0_1_wdata;
  wire ram_w16_l1024_id9_0_1_wenable;
  wire ram_w16_l1024_id9_0_1_enable;
  assign ram_w16_l1024_id9_0_0_addr = 'hx;
  assign ram_w16_l1024_id9_0_0_wdata = 'hx;
  assign ram_w16_l1024_id9_0_0_wenable = 0;
  assign ram_w16_l1024_id9_0_0_enable = 0;
  assign ram_w16_l1024_id9_0_1_addr = 'hx;
  assign ram_w16_l1024_id9_0_1_wdata = 'hx;
  assign ram_w16_l1024_id9_0_1_wenable = 0;
  assign ram_w16_l1024_id9_0_1_enable = 0;

  ram_w16_l1024_id9_0
  inst_ram_w16_l1024_id9_0
  (
    .CLK(CLK),
    .ram_w16_l1024_id9_0_0_addr(ram_w16_l1024_id9_0_0_addr),
    .ram_w16_l1024_id9_0_0_rdata(ram_w16_l1024_id9_0_0_rdata),
    .ram_w16_l1024_id9_0_0_wdata(ram_w16_l1024_id9_0_0_wdata),
    .ram_w16_l1024_id9_0_0_wenable(ram_w16_l1024_id9_0_0_wenable),
    .ram_w16_l1024_id9_0_0_enable(ram_w16_l1024_id9_0_0_enable),
    .ram_w16_l1024_id9_0_1_addr(ram_w16_l1024_id9_0_1_addr),
    .ram_w16_l1024_id9_0_1_rdata(ram_w16_l1024_id9_0_1_rdata),
    .ram_w16_l1024_id9_0_1_wdata(ram_w16_l1024_id9_0_1_wdata),
    .ram_w16_l1024_id9_0_1_wenable(ram_w16_l1024_id9_0_1_wenable),
    .ram_w16_l1024_id9_0_1_enable(ram_w16_l1024_id9_0_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id9_1_0_addr;
  wire [16-1:0] ram_w16_l1024_id9_1_0_rdata;
  wire [16-1:0] ram_w16_l1024_id9_1_0_wdata;
  wire ram_w16_l1024_id9_1_0_wenable;
  wire ram_w16_l1024_id9_1_0_enable;
  wire [9-1:0] ram_w16_l1024_id9_1_1_addr;
  wire [16-1:0] ram_w16_l1024_id9_1_1_rdata;
  wire [16-1:0] ram_w16_l1024_id9_1_1_wdata;
  wire ram_w16_l1024_id9_1_1_wenable;
  wire ram_w16_l1024_id9_1_1_enable;
  assign ram_w16_l1024_id9_1_0_addr = 'hx;
  assign ram_w16_l1024_id9_1_0_wdata = 'hx;
  assign ram_w16_l1024_id9_1_0_wenable = 0;
  assign ram_w16_l1024_id9_1_0_enable = 0;
  assign ram_w16_l1024_id9_1_1_addr = 'hx;
  assign ram_w16_l1024_id9_1_1_wdata = 'hx;
  assign ram_w16_l1024_id9_1_1_wenable = 0;
  assign ram_w16_l1024_id9_1_1_enable = 0;

  ram_w16_l1024_id9_1
  inst_ram_w16_l1024_id9_1
  (
    .CLK(CLK),
    .ram_w16_l1024_id9_1_0_addr(ram_w16_l1024_id9_1_0_addr),
    .ram_w16_l1024_id9_1_0_rdata(ram_w16_l1024_id9_1_0_rdata),
    .ram_w16_l1024_id9_1_0_wdata(ram_w16_l1024_id9_1_0_wdata),
    .ram_w16_l1024_id9_1_0_wenable(ram_w16_l1024_id9_1_0_wenable),
    .ram_w16_l1024_id9_1_0_enable(ram_w16_l1024_id9_1_0_enable),
    .ram_w16_l1024_id9_1_1_addr(ram_w16_l1024_id9_1_1_addr),
    .ram_w16_l1024_id9_1_1_rdata(ram_w16_l1024_id9_1_1_rdata),
    .ram_w16_l1024_id9_1_1_wdata(ram_w16_l1024_id9_1_1_wdata),
    .ram_w16_l1024_id9_1_1_wenable(ram_w16_l1024_id9_1_1_wenable),
    .ram_w16_l1024_id9_1_1_enable(ram_w16_l1024_id9_1_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id10_0_0_addr;
  wire [16-1:0] ram_w16_l1024_id10_0_0_rdata;
  wire [16-1:0] ram_w16_l1024_id10_0_0_wdata;
  wire ram_w16_l1024_id10_0_0_wenable;
  wire ram_w16_l1024_id10_0_0_enable;
  wire [9-1:0] ram_w16_l1024_id10_0_1_addr;
  wire [16-1:0] ram_w16_l1024_id10_0_1_rdata;
  wire [16-1:0] ram_w16_l1024_id10_0_1_wdata;
  wire ram_w16_l1024_id10_0_1_wenable;
  wire ram_w16_l1024_id10_0_1_enable;
  assign ram_w16_l1024_id10_0_0_addr = 'hx;
  assign ram_w16_l1024_id10_0_0_wdata = 'hx;
  assign ram_w16_l1024_id10_0_0_wenable = 0;
  assign ram_w16_l1024_id10_0_0_enable = 0;
  assign ram_w16_l1024_id10_0_1_addr = 'hx;
  assign ram_w16_l1024_id10_0_1_wdata = 'hx;
  assign ram_w16_l1024_id10_0_1_wenable = 0;
  assign ram_w16_l1024_id10_0_1_enable = 0;

  ram_w16_l1024_id10_0
  inst_ram_w16_l1024_id10_0
  (
    .CLK(CLK),
    .ram_w16_l1024_id10_0_0_addr(ram_w16_l1024_id10_0_0_addr),
    .ram_w16_l1024_id10_0_0_rdata(ram_w16_l1024_id10_0_0_rdata),
    .ram_w16_l1024_id10_0_0_wdata(ram_w16_l1024_id10_0_0_wdata),
    .ram_w16_l1024_id10_0_0_wenable(ram_w16_l1024_id10_0_0_wenable),
    .ram_w16_l1024_id10_0_0_enable(ram_w16_l1024_id10_0_0_enable),
    .ram_w16_l1024_id10_0_1_addr(ram_w16_l1024_id10_0_1_addr),
    .ram_w16_l1024_id10_0_1_rdata(ram_w16_l1024_id10_0_1_rdata),
    .ram_w16_l1024_id10_0_1_wdata(ram_w16_l1024_id10_0_1_wdata),
    .ram_w16_l1024_id10_0_1_wenable(ram_w16_l1024_id10_0_1_wenable),
    .ram_w16_l1024_id10_0_1_enable(ram_w16_l1024_id10_0_1_enable)
  );

  wire [9-1:0] ram_w16_l1024_id10_1_0_addr;
  wire [16-1:0] ram_w16_l1024_id10_1_0_rdata;
  wire [16-1:0] ram_w16_l1024_id10_1_0_wdata;
  wire ram_w16_l1024_id10_1_0_wenable;
  wire ram_w16_l1024_id10_1_0_enable;
  wire [9-1:0] ram_w16_l1024_id10_1_1_addr;
  wire [16-1:0] ram_w16_l1024_id10_1_1_rdata;
  wire [16-1:0] ram_w16_l1024_id10_1_1_wdata;
  wire ram_w16_l1024_id10_1_1_wenable;
  wire ram_w16_l1024_id10_1_1_enable;
  assign ram_w16_l1024_id10_1_0_addr = 'hx;
  assign ram_w16_l1024_id10_1_0_wdata = 'hx;
  assign ram_w16_l1024_id10_1_0_wenable = 0;
  assign ram_w16_l1024_id10_1_0_enable = 0;
  assign ram_w16_l1024_id10_1_1_addr = 'hx;
  assign ram_w16_l1024_id10_1_1_wdata = 'hx;
  assign ram_w16_l1024_id10_1_1_wenable = 0;
  assign ram_w16_l1024_id10_1_1_enable = 0;

  ram_w16_l1024_id10_1
  inst_ram_w16_l1024_id10_1
  (
    .CLK(CLK),
    .ram_w16_l1024_id10_1_0_addr(ram_w16_l1024_id10_1_0_addr),
    .ram_w16_l1024_id10_1_0_rdata(ram_w16_l1024_id10_1_0_rdata),
    .ram_w16_l1024_id10_1_0_wdata(ram_w16_l1024_id10_1_0_wdata),
    .ram_w16_l1024_id10_1_0_wenable(ram_w16_l1024_id10_1_0_wenable),
    .ram_w16_l1024_id10_1_0_enable(ram_w16_l1024_id10_1_0_enable),
    .ram_w16_l1024_id10_1_1_addr(ram_w16_l1024_id10_1_1_addr),
    .ram_w16_l1024_id10_1_1_rdata(ram_w16_l1024_id10_1_1_rdata),
    .ram_w16_l1024_id10_1_1_wdata(ram_w16_l1024_id10_1_1_wdata),
    .ram_w16_l1024_id10_1_1_wenable(ram_w16_l1024_id10_1_1_wenable),
    .ram_w16_l1024_id10_1_1_enable(ram_w16_l1024_id10_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id0_0_0_addr;
  wire [16-1:0] ram_w16_l512_id0_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id0_0_0_wdata;
  wire ram_w16_l512_id0_0_0_wenable;
  wire ram_w16_l512_id0_0_0_enable;
  wire [8-1:0] ram_w16_l512_id0_0_1_addr;
  wire [16-1:0] ram_w16_l512_id0_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id0_0_1_wdata;
  wire ram_w16_l512_id0_0_1_wenable;
  wire ram_w16_l512_id0_0_1_enable;
  assign ram_w16_l512_id0_0_1_wdata = 'hx;
  assign ram_w16_l512_id0_0_1_wenable = 0;

  ram_w16_l512_id0_0
  inst_ram_w16_l512_id0_0
  (
    .CLK(CLK),
    .ram_w16_l512_id0_0_0_addr(ram_w16_l512_id0_0_0_addr),
    .ram_w16_l512_id0_0_0_rdata(ram_w16_l512_id0_0_0_rdata),
    .ram_w16_l512_id0_0_0_wdata(ram_w16_l512_id0_0_0_wdata),
    .ram_w16_l512_id0_0_0_wenable(ram_w16_l512_id0_0_0_wenable),
    .ram_w16_l512_id0_0_0_enable(ram_w16_l512_id0_0_0_enable),
    .ram_w16_l512_id0_0_1_addr(ram_w16_l512_id0_0_1_addr),
    .ram_w16_l512_id0_0_1_rdata(ram_w16_l512_id0_0_1_rdata),
    .ram_w16_l512_id0_0_1_wdata(ram_w16_l512_id0_0_1_wdata),
    .ram_w16_l512_id0_0_1_wenable(ram_w16_l512_id0_0_1_wenable),
    .ram_w16_l512_id0_0_1_enable(ram_w16_l512_id0_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id0_1_0_addr;
  wire [16-1:0] ram_w16_l512_id0_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id0_1_0_wdata;
  wire ram_w16_l512_id0_1_0_wenable;
  wire ram_w16_l512_id0_1_0_enable;
  wire [8-1:0] ram_w16_l512_id0_1_1_addr;
  wire [16-1:0] ram_w16_l512_id0_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id0_1_1_wdata;
  wire ram_w16_l512_id0_1_1_wenable;
  wire ram_w16_l512_id0_1_1_enable;
  assign ram_w16_l512_id0_1_1_wdata = 'hx;
  assign ram_w16_l512_id0_1_1_wenable = 0;

  ram_w16_l512_id0_1
  inst_ram_w16_l512_id0_1
  (
    .CLK(CLK),
    .ram_w16_l512_id0_1_0_addr(ram_w16_l512_id0_1_0_addr),
    .ram_w16_l512_id0_1_0_rdata(ram_w16_l512_id0_1_0_rdata),
    .ram_w16_l512_id0_1_0_wdata(ram_w16_l512_id0_1_0_wdata),
    .ram_w16_l512_id0_1_0_wenable(ram_w16_l512_id0_1_0_wenable),
    .ram_w16_l512_id0_1_0_enable(ram_w16_l512_id0_1_0_enable),
    .ram_w16_l512_id0_1_1_addr(ram_w16_l512_id0_1_1_addr),
    .ram_w16_l512_id0_1_1_rdata(ram_w16_l512_id0_1_1_rdata),
    .ram_w16_l512_id0_1_1_wdata(ram_w16_l512_id0_1_1_wdata),
    .ram_w16_l512_id0_1_1_wenable(ram_w16_l512_id0_1_1_wenable),
    .ram_w16_l512_id0_1_1_enable(ram_w16_l512_id0_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id1_0_0_addr;
  wire [16-1:0] ram_w16_l512_id1_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id1_0_0_wdata;
  wire ram_w16_l512_id1_0_0_wenable;
  wire ram_w16_l512_id1_0_0_enable;
  wire [8-1:0] ram_w16_l512_id1_0_1_addr;
  wire [16-1:0] ram_w16_l512_id1_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id1_0_1_wdata;
  wire ram_w16_l512_id1_0_1_wenable;
  wire ram_w16_l512_id1_0_1_enable;
  assign ram_w16_l512_id1_0_0_wdata = 'hx;
  assign ram_w16_l512_id1_0_0_wenable = 0;

  ram_w16_l512_id1_0
  inst_ram_w16_l512_id1_0
  (
    .CLK(CLK),
    .ram_w16_l512_id1_0_0_addr(ram_w16_l512_id1_0_0_addr),
    .ram_w16_l512_id1_0_0_rdata(ram_w16_l512_id1_0_0_rdata),
    .ram_w16_l512_id1_0_0_wdata(ram_w16_l512_id1_0_0_wdata),
    .ram_w16_l512_id1_0_0_wenable(ram_w16_l512_id1_0_0_wenable),
    .ram_w16_l512_id1_0_0_enable(ram_w16_l512_id1_0_0_enable),
    .ram_w16_l512_id1_0_1_addr(ram_w16_l512_id1_0_1_addr),
    .ram_w16_l512_id1_0_1_rdata(ram_w16_l512_id1_0_1_rdata),
    .ram_w16_l512_id1_0_1_wdata(ram_w16_l512_id1_0_1_wdata),
    .ram_w16_l512_id1_0_1_wenable(ram_w16_l512_id1_0_1_wenable),
    .ram_w16_l512_id1_0_1_enable(ram_w16_l512_id1_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id1_1_0_addr;
  wire [16-1:0] ram_w16_l512_id1_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id1_1_0_wdata;
  wire ram_w16_l512_id1_1_0_wenable;
  wire ram_w16_l512_id1_1_0_enable;
  wire [8-1:0] ram_w16_l512_id1_1_1_addr;
  wire [16-1:0] ram_w16_l512_id1_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id1_1_1_wdata;
  wire ram_w16_l512_id1_1_1_wenable;
  wire ram_w16_l512_id1_1_1_enable;
  assign ram_w16_l512_id1_1_0_wdata = 'hx;
  assign ram_w16_l512_id1_1_0_wenable = 0;

  ram_w16_l512_id1_1
  inst_ram_w16_l512_id1_1
  (
    .CLK(CLK),
    .ram_w16_l512_id1_1_0_addr(ram_w16_l512_id1_1_0_addr),
    .ram_w16_l512_id1_1_0_rdata(ram_w16_l512_id1_1_0_rdata),
    .ram_w16_l512_id1_1_0_wdata(ram_w16_l512_id1_1_0_wdata),
    .ram_w16_l512_id1_1_0_wenable(ram_w16_l512_id1_1_0_wenable),
    .ram_w16_l512_id1_1_0_enable(ram_w16_l512_id1_1_0_enable),
    .ram_w16_l512_id1_1_1_addr(ram_w16_l512_id1_1_1_addr),
    .ram_w16_l512_id1_1_1_rdata(ram_w16_l512_id1_1_1_rdata),
    .ram_w16_l512_id1_1_1_wdata(ram_w16_l512_id1_1_1_wdata),
    .ram_w16_l512_id1_1_1_wenable(ram_w16_l512_id1_1_1_wenable),
    .ram_w16_l512_id1_1_1_enable(ram_w16_l512_id1_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id2_0_0_addr;
  wire [16-1:0] ram_w16_l512_id2_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id2_0_0_wdata;
  wire ram_w16_l512_id2_0_0_wenable;
  wire ram_w16_l512_id2_0_0_enable;
  wire [8-1:0] ram_w16_l512_id2_0_1_addr;
  wire [16-1:0] ram_w16_l512_id2_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id2_0_1_wdata;
  wire ram_w16_l512_id2_0_1_wenable;
  wire ram_w16_l512_id2_0_1_enable;
  assign ram_w16_l512_id2_0_0_wdata = 'hx;
  assign ram_w16_l512_id2_0_0_wenable = 0;

  ram_w16_l512_id2_0
  inst_ram_w16_l512_id2_0
  (
    .CLK(CLK),
    .ram_w16_l512_id2_0_0_addr(ram_w16_l512_id2_0_0_addr),
    .ram_w16_l512_id2_0_0_rdata(ram_w16_l512_id2_0_0_rdata),
    .ram_w16_l512_id2_0_0_wdata(ram_w16_l512_id2_0_0_wdata),
    .ram_w16_l512_id2_0_0_wenable(ram_w16_l512_id2_0_0_wenable),
    .ram_w16_l512_id2_0_0_enable(ram_w16_l512_id2_0_0_enable),
    .ram_w16_l512_id2_0_1_addr(ram_w16_l512_id2_0_1_addr),
    .ram_w16_l512_id2_0_1_rdata(ram_w16_l512_id2_0_1_rdata),
    .ram_w16_l512_id2_0_1_wdata(ram_w16_l512_id2_0_1_wdata),
    .ram_w16_l512_id2_0_1_wenable(ram_w16_l512_id2_0_1_wenable),
    .ram_w16_l512_id2_0_1_enable(ram_w16_l512_id2_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id2_1_0_addr;
  wire [16-1:0] ram_w16_l512_id2_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id2_1_0_wdata;
  wire ram_w16_l512_id2_1_0_wenable;
  wire ram_w16_l512_id2_1_0_enable;
  wire [8-1:0] ram_w16_l512_id2_1_1_addr;
  wire [16-1:0] ram_w16_l512_id2_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id2_1_1_wdata;
  wire ram_w16_l512_id2_1_1_wenable;
  wire ram_w16_l512_id2_1_1_enable;
  assign ram_w16_l512_id2_1_0_wdata = 'hx;
  assign ram_w16_l512_id2_1_0_wenable = 0;

  ram_w16_l512_id2_1
  inst_ram_w16_l512_id2_1
  (
    .CLK(CLK),
    .ram_w16_l512_id2_1_0_addr(ram_w16_l512_id2_1_0_addr),
    .ram_w16_l512_id2_1_0_rdata(ram_w16_l512_id2_1_0_rdata),
    .ram_w16_l512_id2_1_0_wdata(ram_w16_l512_id2_1_0_wdata),
    .ram_w16_l512_id2_1_0_wenable(ram_w16_l512_id2_1_0_wenable),
    .ram_w16_l512_id2_1_0_enable(ram_w16_l512_id2_1_0_enable),
    .ram_w16_l512_id2_1_1_addr(ram_w16_l512_id2_1_1_addr),
    .ram_w16_l512_id2_1_1_rdata(ram_w16_l512_id2_1_1_rdata),
    .ram_w16_l512_id2_1_1_wdata(ram_w16_l512_id2_1_1_wdata),
    .ram_w16_l512_id2_1_1_wenable(ram_w16_l512_id2_1_1_wenable),
    .ram_w16_l512_id2_1_1_enable(ram_w16_l512_id2_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id3_0_0_addr;
  wire [16-1:0] ram_w16_l512_id3_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id3_0_0_wdata;
  wire ram_w16_l512_id3_0_0_wenable;
  wire ram_w16_l512_id3_0_0_enable;
  wire [8-1:0] ram_w16_l512_id3_0_1_addr;
  wire [16-1:0] ram_w16_l512_id3_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id3_0_1_wdata;
  wire ram_w16_l512_id3_0_1_wenable;
  wire ram_w16_l512_id3_0_1_enable;
  assign ram_w16_l512_id3_0_0_wdata = 'hx;
  assign ram_w16_l512_id3_0_0_wenable = 0;

  ram_w16_l512_id3_0
  inst_ram_w16_l512_id3_0
  (
    .CLK(CLK),
    .ram_w16_l512_id3_0_0_addr(ram_w16_l512_id3_0_0_addr),
    .ram_w16_l512_id3_0_0_rdata(ram_w16_l512_id3_0_0_rdata),
    .ram_w16_l512_id3_0_0_wdata(ram_w16_l512_id3_0_0_wdata),
    .ram_w16_l512_id3_0_0_wenable(ram_w16_l512_id3_0_0_wenable),
    .ram_w16_l512_id3_0_0_enable(ram_w16_l512_id3_0_0_enable),
    .ram_w16_l512_id3_0_1_addr(ram_w16_l512_id3_0_1_addr),
    .ram_w16_l512_id3_0_1_rdata(ram_w16_l512_id3_0_1_rdata),
    .ram_w16_l512_id3_0_1_wdata(ram_w16_l512_id3_0_1_wdata),
    .ram_w16_l512_id3_0_1_wenable(ram_w16_l512_id3_0_1_wenable),
    .ram_w16_l512_id3_0_1_enable(ram_w16_l512_id3_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id3_1_0_addr;
  wire [16-1:0] ram_w16_l512_id3_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id3_1_0_wdata;
  wire ram_w16_l512_id3_1_0_wenable;
  wire ram_w16_l512_id3_1_0_enable;
  wire [8-1:0] ram_w16_l512_id3_1_1_addr;
  wire [16-1:0] ram_w16_l512_id3_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id3_1_1_wdata;
  wire ram_w16_l512_id3_1_1_wenable;
  wire ram_w16_l512_id3_1_1_enable;
  assign ram_w16_l512_id3_1_0_wdata = 'hx;
  assign ram_w16_l512_id3_1_0_wenable = 0;

  ram_w16_l512_id3_1
  inst_ram_w16_l512_id3_1
  (
    .CLK(CLK),
    .ram_w16_l512_id3_1_0_addr(ram_w16_l512_id3_1_0_addr),
    .ram_w16_l512_id3_1_0_rdata(ram_w16_l512_id3_1_0_rdata),
    .ram_w16_l512_id3_1_0_wdata(ram_w16_l512_id3_1_0_wdata),
    .ram_w16_l512_id3_1_0_wenable(ram_w16_l512_id3_1_0_wenable),
    .ram_w16_l512_id3_1_0_enable(ram_w16_l512_id3_1_0_enable),
    .ram_w16_l512_id3_1_1_addr(ram_w16_l512_id3_1_1_addr),
    .ram_w16_l512_id3_1_1_rdata(ram_w16_l512_id3_1_1_rdata),
    .ram_w16_l512_id3_1_1_wdata(ram_w16_l512_id3_1_1_wdata),
    .ram_w16_l512_id3_1_1_wenable(ram_w16_l512_id3_1_1_wenable),
    .ram_w16_l512_id3_1_1_enable(ram_w16_l512_id3_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id4_0_0_addr;
  wire [16-1:0] ram_w16_l512_id4_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id4_0_0_wdata;
  wire ram_w16_l512_id4_0_0_wenable;
  wire ram_w16_l512_id4_0_0_enable;
  wire [8-1:0] ram_w16_l512_id4_0_1_addr;
  wire [16-1:0] ram_w16_l512_id4_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id4_0_1_wdata;
  wire ram_w16_l512_id4_0_1_wenable;
  wire ram_w16_l512_id4_0_1_enable;
  assign ram_w16_l512_id4_0_0_wdata = 'hx;
  assign ram_w16_l512_id4_0_0_wenable = 0;

  ram_w16_l512_id4_0
  inst_ram_w16_l512_id4_0
  (
    .CLK(CLK),
    .ram_w16_l512_id4_0_0_addr(ram_w16_l512_id4_0_0_addr),
    .ram_w16_l512_id4_0_0_rdata(ram_w16_l512_id4_0_0_rdata),
    .ram_w16_l512_id4_0_0_wdata(ram_w16_l512_id4_0_0_wdata),
    .ram_w16_l512_id4_0_0_wenable(ram_w16_l512_id4_0_0_wenable),
    .ram_w16_l512_id4_0_0_enable(ram_w16_l512_id4_0_0_enable),
    .ram_w16_l512_id4_0_1_addr(ram_w16_l512_id4_0_1_addr),
    .ram_w16_l512_id4_0_1_rdata(ram_w16_l512_id4_0_1_rdata),
    .ram_w16_l512_id4_0_1_wdata(ram_w16_l512_id4_0_1_wdata),
    .ram_w16_l512_id4_0_1_wenable(ram_w16_l512_id4_0_1_wenable),
    .ram_w16_l512_id4_0_1_enable(ram_w16_l512_id4_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id4_1_0_addr;
  wire [16-1:0] ram_w16_l512_id4_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id4_1_0_wdata;
  wire ram_w16_l512_id4_1_0_wenable;
  wire ram_w16_l512_id4_1_0_enable;
  wire [8-1:0] ram_w16_l512_id4_1_1_addr;
  wire [16-1:0] ram_w16_l512_id4_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id4_1_1_wdata;
  wire ram_w16_l512_id4_1_1_wenable;
  wire ram_w16_l512_id4_1_1_enable;
  assign ram_w16_l512_id4_1_0_wdata = 'hx;
  assign ram_w16_l512_id4_1_0_wenable = 0;

  ram_w16_l512_id4_1
  inst_ram_w16_l512_id4_1
  (
    .CLK(CLK),
    .ram_w16_l512_id4_1_0_addr(ram_w16_l512_id4_1_0_addr),
    .ram_w16_l512_id4_1_0_rdata(ram_w16_l512_id4_1_0_rdata),
    .ram_w16_l512_id4_1_0_wdata(ram_w16_l512_id4_1_0_wdata),
    .ram_w16_l512_id4_1_0_wenable(ram_w16_l512_id4_1_0_wenable),
    .ram_w16_l512_id4_1_0_enable(ram_w16_l512_id4_1_0_enable),
    .ram_w16_l512_id4_1_1_addr(ram_w16_l512_id4_1_1_addr),
    .ram_w16_l512_id4_1_1_rdata(ram_w16_l512_id4_1_1_rdata),
    .ram_w16_l512_id4_1_1_wdata(ram_w16_l512_id4_1_1_wdata),
    .ram_w16_l512_id4_1_1_wenable(ram_w16_l512_id4_1_1_wenable),
    .ram_w16_l512_id4_1_1_enable(ram_w16_l512_id4_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id5_0_0_addr;
  wire [16-1:0] ram_w16_l512_id5_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id5_0_0_wdata;
  wire ram_w16_l512_id5_0_0_wenable;
  wire ram_w16_l512_id5_0_0_enable;
  wire [8-1:0] ram_w16_l512_id5_0_1_addr;
  wire [16-1:0] ram_w16_l512_id5_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id5_0_1_wdata;
  wire ram_w16_l512_id5_0_1_wenable;
  wire ram_w16_l512_id5_0_1_enable;
  assign ram_w16_l512_id5_0_0_wdata = 'hx;
  assign ram_w16_l512_id5_0_0_wenable = 0;

  ram_w16_l512_id5_0
  inst_ram_w16_l512_id5_0
  (
    .CLK(CLK),
    .ram_w16_l512_id5_0_0_addr(ram_w16_l512_id5_0_0_addr),
    .ram_w16_l512_id5_0_0_rdata(ram_w16_l512_id5_0_0_rdata),
    .ram_w16_l512_id5_0_0_wdata(ram_w16_l512_id5_0_0_wdata),
    .ram_w16_l512_id5_0_0_wenable(ram_w16_l512_id5_0_0_wenable),
    .ram_w16_l512_id5_0_0_enable(ram_w16_l512_id5_0_0_enable),
    .ram_w16_l512_id5_0_1_addr(ram_w16_l512_id5_0_1_addr),
    .ram_w16_l512_id5_0_1_rdata(ram_w16_l512_id5_0_1_rdata),
    .ram_w16_l512_id5_0_1_wdata(ram_w16_l512_id5_0_1_wdata),
    .ram_w16_l512_id5_0_1_wenable(ram_w16_l512_id5_0_1_wenable),
    .ram_w16_l512_id5_0_1_enable(ram_w16_l512_id5_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id5_1_0_addr;
  wire [16-1:0] ram_w16_l512_id5_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id5_1_0_wdata;
  wire ram_w16_l512_id5_1_0_wenable;
  wire ram_w16_l512_id5_1_0_enable;
  wire [8-1:0] ram_w16_l512_id5_1_1_addr;
  wire [16-1:0] ram_w16_l512_id5_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id5_1_1_wdata;
  wire ram_w16_l512_id5_1_1_wenable;
  wire ram_w16_l512_id5_1_1_enable;
  assign ram_w16_l512_id5_1_0_wdata = 'hx;
  assign ram_w16_l512_id5_1_0_wenable = 0;

  ram_w16_l512_id5_1
  inst_ram_w16_l512_id5_1
  (
    .CLK(CLK),
    .ram_w16_l512_id5_1_0_addr(ram_w16_l512_id5_1_0_addr),
    .ram_w16_l512_id5_1_0_rdata(ram_w16_l512_id5_1_0_rdata),
    .ram_w16_l512_id5_1_0_wdata(ram_w16_l512_id5_1_0_wdata),
    .ram_w16_l512_id5_1_0_wenable(ram_w16_l512_id5_1_0_wenable),
    .ram_w16_l512_id5_1_0_enable(ram_w16_l512_id5_1_0_enable),
    .ram_w16_l512_id5_1_1_addr(ram_w16_l512_id5_1_1_addr),
    .ram_w16_l512_id5_1_1_rdata(ram_w16_l512_id5_1_1_rdata),
    .ram_w16_l512_id5_1_1_wdata(ram_w16_l512_id5_1_1_wdata),
    .ram_w16_l512_id5_1_1_wenable(ram_w16_l512_id5_1_1_wenable),
    .ram_w16_l512_id5_1_1_enable(ram_w16_l512_id5_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id6_0_0_addr;
  wire [16-1:0] ram_w16_l512_id6_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id6_0_0_wdata;
  wire ram_w16_l512_id6_0_0_wenable;
  wire ram_w16_l512_id6_0_0_enable;
  wire [8-1:0] ram_w16_l512_id6_0_1_addr;
  wire [16-1:0] ram_w16_l512_id6_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id6_0_1_wdata;
  wire ram_w16_l512_id6_0_1_wenable;
  wire ram_w16_l512_id6_0_1_enable;
  assign ram_w16_l512_id6_0_0_wdata = 'hx;
  assign ram_w16_l512_id6_0_0_wenable = 0;

  ram_w16_l512_id6_0
  inst_ram_w16_l512_id6_0
  (
    .CLK(CLK),
    .ram_w16_l512_id6_0_0_addr(ram_w16_l512_id6_0_0_addr),
    .ram_w16_l512_id6_0_0_rdata(ram_w16_l512_id6_0_0_rdata),
    .ram_w16_l512_id6_0_0_wdata(ram_w16_l512_id6_0_0_wdata),
    .ram_w16_l512_id6_0_0_wenable(ram_w16_l512_id6_0_0_wenable),
    .ram_w16_l512_id6_0_0_enable(ram_w16_l512_id6_0_0_enable),
    .ram_w16_l512_id6_0_1_addr(ram_w16_l512_id6_0_1_addr),
    .ram_w16_l512_id6_0_1_rdata(ram_w16_l512_id6_0_1_rdata),
    .ram_w16_l512_id6_0_1_wdata(ram_w16_l512_id6_0_1_wdata),
    .ram_w16_l512_id6_0_1_wenable(ram_w16_l512_id6_0_1_wenable),
    .ram_w16_l512_id6_0_1_enable(ram_w16_l512_id6_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id6_1_0_addr;
  wire [16-1:0] ram_w16_l512_id6_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id6_1_0_wdata;
  wire ram_w16_l512_id6_1_0_wenable;
  wire ram_w16_l512_id6_1_0_enable;
  wire [8-1:0] ram_w16_l512_id6_1_1_addr;
  wire [16-1:0] ram_w16_l512_id6_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id6_1_1_wdata;
  wire ram_w16_l512_id6_1_1_wenable;
  wire ram_w16_l512_id6_1_1_enable;
  assign ram_w16_l512_id6_1_0_wdata = 'hx;
  assign ram_w16_l512_id6_1_0_wenable = 0;

  ram_w16_l512_id6_1
  inst_ram_w16_l512_id6_1
  (
    .CLK(CLK),
    .ram_w16_l512_id6_1_0_addr(ram_w16_l512_id6_1_0_addr),
    .ram_w16_l512_id6_1_0_rdata(ram_w16_l512_id6_1_0_rdata),
    .ram_w16_l512_id6_1_0_wdata(ram_w16_l512_id6_1_0_wdata),
    .ram_w16_l512_id6_1_0_wenable(ram_w16_l512_id6_1_0_wenable),
    .ram_w16_l512_id6_1_0_enable(ram_w16_l512_id6_1_0_enable),
    .ram_w16_l512_id6_1_1_addr(ram_w16_l512_id6_1_1_addr),
    .ram_w16_l512_id6_1_1_rdata(ram_w16_l512_id6_1_1_rdata),
    .ram_w16_l512_id6_1_1_wdata(ram_w16_l512_id6_1_1_wdata),
    .ram_w16_l512_id6_1_1_wenable(ram_w16_l512_id6_1_1_wenable),
    .ram_w16_l512_id6_1_1_enable(ram_w16_l512_id6_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id7_0_0_addr;
  wire [16-1:0] ram_w16_l512_id7_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id7_0_0_wdata;
  wire ram_w16_l512_id7_0_0_wenable;
  wire ram_w16_l512_id7_0_0_enable;
  wire [8-1:0] ram_w16_l512_id7_0_1_addr;
  wire [16-1:0] ram_w16_l512_id7_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id7_0_1_wdata;
  wire ram_w16_l512_id7_0_1_wenable;
  wire ram_w16_l512_id7_0_1_enable;
  assign ram_w16_l512_id7_0_0_wdata = 'hx;
  assign ram_w16_l512_id7_0_0_wenable = 0;

  ram_w16_l512_id7_0
  inst_ram_w16_l512_id7_0
  (
    .CLK(CLK),
    .ram_w16_l512_id7_0_0_addr(ram_w16_l512_id7_0_0_addr),
    .ram_w16_l512_id7_0_0_rdata(ram_w16_l512_id7_0_0_rdata),
    .ram_w16_l512_id7_0_0_wdata(ram_w16_l512_id7_0_0_wdata),
    .ram_w16_l512_id7_0_0_wenable(ram_w16_l512_id7_0_0_wenable),
    .ram_w16_l512_id7_0_0_enable(ram_w16_l512_id7_0_0_enable),
    .ram_w16_l512_id7_0_1_addr(ram_w16_l512_id7_0_1_addr),
    .ram_w16_l512_id7_0_1_rdata(ram_w16_l512_id7_0_1_rdata),
    .ram_w16_l512_id7_0_1_wdata(ram_w16_l512_id7_0_1_wdata),
    .ram_w16_l512_id7_0_1_wenable(ram_w16_l512_id7_0_1_wenable),
    .ram_w16_l512_id7_0_1_enable(ram_w16_l512_id7_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id7_1_0_addr;
  wire [16-1:0] ram_w16_l512_id7_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id7_1_0_wdata;
  wire ram_w16_l512_id7_1_0_wenable;
  wire ram_w16_l512_id7_1_0_enable;
  wire [8-1:0] ram_w16_l512_id7_1_1_addr;
  wire [16-1:0] ram_w16_l512_id7_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id7_1_1_wdata;
  wire ram_w16_l512_id7_1_1_wenable;
  wire ram_w16_l512_id7_1_1_enable;
  assign ram_w16_l512_id7_1_0_wdata = 'hx;
  assign ram_w16_l512_id7_1_0_wenable = 0;

  ram_w16_l512_id7_1
  inst_ram_w16_l512_id7_1
  (
    .CLK(CLK),
    .ram_w16_l512_id7_1_0_addr(ram_w16_l512_id7_1_0_addr),
    .ram_w16_l512_id7_1_0_rdata(ram_w16_l512_id7_1_0_rdata),
    .ram_w16_l512_id7_1_0_wdata(ram_w16_l512_id7_1_0_wdata),
    .ram_w16_l512_id7_1_0_wenable(ram_w16_l512_id7_1_0_wenable),
    .ram_w16_l512_id7_1_0_enable(ram_w16_l512_id7_1_0_enable),
    .ram_w16_l512_id7_1_1_addr(ram_w16_l512_id7_1_1_addr),
    .ram_w16_l512_id7_1_1_rdata(ram_w16_l512_id7_1_1_rdata),
    .ram_w16_l512_id7_1_1_wdata(ram_w16_l512_id7_1_1_wdata),
    .ram_w16_l512_id7_1_1_wenable(ram_w16_l512_id7_1_1_wenable),
    .ram_w16_l512_id7_1_1_enable(ram_w16_l512_id7_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id8_0_0_addr;
  wire [16-1:0] ram_w16_l512_id8_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id8_0_0_wdata;
  wire ram_w16_l512_id8_0_0_wenable;
  wire ram_w16_l512_id8_0_0_enable;
  wire [8-1:0] ram_w16_l512_id8_0_1_addr;
  wire [16-1:0] ram_w16_l512_id8_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id8_0_1_wdata;
  wire ram_w16_l512_id8_0_1_wenable;
  wire ram_w16_l512_id8_0_1_enable;
  assign ram_w16_l512_id8_0_0_wdata = 'hx;
  assign ram_w16_l512_id8_0_0_wenable = 0;

  ram_w16_l512_id8_0
  inst_ram_w16_l512_id8_0
  (
    .CLK(CLK),
    .ram_w16_l512_id8_0_0_addr(ram_w16_l512_id8_0_0_addr),
    .ram_w16_l512_id8_0_0_rdata(ram_w16_l512_id8_0_0_rdata),
    .ram_w16_l512_id8_0_0_wdata(ram_w16_l512_id8_0_0_wdata),
    .ram_w16_l512_id8_0_0_wenable(ram_w16_l512_id8_0_0_wenable),
    .ram_w16_l512_id8_0_0_enable(ram_w16_l512_id8_0_0_enable),
    .ram_w16_l512_id8_0_1_addr(ram_w16_l512_id8_0_1_addr),
    .ram_w16_l512_id8_0_1_rdata(ram_w16_l512_id8_0_1_rdata),
    .ram_w16_l512_id8_0_1_wdata(ram_w16_l512_id8_0_1_wdata),
    .ram_w16_l512_id8_0_1_wenable(ram_w16_l512_id8_0_1_wenable),
    .ram_w16_l512_id8_0_1_enable(ram_w16_l512_id8_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id8_1_0_addr;
  wire [16-1:0] ram_w16_l512_id8_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id8_1_0_wdata;
  wire ram_w16_l512_id8_1_0_wenable;
  wire ram_w16_l512_id8_1_0_enable;
  wire [8-1:0] ram_w16_l512_id8_1_1_addr;
  wire [16-1:0] ram_w16_l512_id8_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id8_1_1_wdata;
  wire ram_w16_l512_id8_1_1_wenable;
  wire ram_w16_l512_id8_1_1_enable;
  assign ram_w16_l512_id8_1_0_wdata = 'hx;
  assign ram_w16_l512_id8_1_0_wenable = 0;

  ram_w16_l512_id8_1
  inst_ram_w16_l512_id8_1
  (
    .CLK(CLK),
    .ram_w16_l512_id8_1_0_addr(ram_w16_l512_id8_1_0_addr),
    .ram_w16_l512_id8_1_0_rdata(ram_w16_l512_id8_1_0_rdata),
    .ram_w16_l512_id8_1_0_wdata(ram_w16_l512_id8_1_0_wdata),
    .ram_w16_l512_id8_1_0_wenable(ram_w16_l512_id8_1_0_wenable),
    .ram_w16_l512_id8_1_0_enable(ram_w16_l512_id8_1_0_enable),
    .ram_w16_l512_id8_1_1_addr(ram_w16_l512_id8_1_1_addr),
    .ram_w16_l512_id8_1_1_rdata(ram_w16_l512_id8_1_1_rdata),
    .ram_w16_l512_id8_1_1_wdata(ram_w16_l512_id8_1_1_wdata),
    .ram_w16_l512_id8_1_1_wenable(ram_w16_l512_id8_1_1_wenable),
    .ram_w16_l512_id8_1_1_enable(ram_w16_l512_id8_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id9_0_0_addr;
  wire [16-1:0] ram_w16_l512_id9_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id9_0_0_wdata;
  wire ram_w16_l512_id9_0_0_wenable;
  wire ram_w16_l512_id9_0_0_enable;
  wire [8-1:0] ram_w16_l512_id9_0_1_addr;
  wire [16-1:0] ram_w16_l512_id9_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id9_0_1_wdata;
  wire ram_w16_l512_id9_0_1_wenable;
  wire ram_w16_l512_id9_0_1_enable;
  assign ram_w16_l512_id9_0_0_wdata = 'hx;
  assign ram_w16_l512_id9_0_0_wenable = 0;

  ram_w16_l512_id9_0
  inst_ram_w16_l512_id9_0
  (
    .CLK(CLK),
    .ram_w16_l512_id9_0_0_addr(ram_w16_l512_id9_0_0_addr),
    .ram_w16_l512_id9_0_0_rdata(ram_w16_l512_id9_0_0_rdata),
    .ram_w16_l512_id9_0_0_wdata(ram_w16_l512_id9_0_0_wdata),
    .ram_w16_l512_id9_0_0_wenable(ram_w16_l512_id9_0_0_wenable),
    .ram_w16_l512_id9_0_0_enable(ram_w16_l512_id9_0_0_enable),
    .ram_w16_l512_id9_0_1_addr(ram_w16_l512_id9_0_1_addr),
    .ram_w16_l512_id9_0_1_rdata(ram_w16_l512_id9_0_1_rdata),
    .ram_w16_l512_id9_0_1_wdata(ram_w16_l512_id9_0_1_wdata),
    .ram_w16_l512_id9_0_1_wenable(ram_w16_l512_id9_0_1_wenable),
    .ram_w16_l512_id9_0_1_enable(ram_w16_l512_id9_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id9_1_0_addr;
  wire [16-1:0] ram_w16_l512_id9_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id9_1_0_wdata;
  wire ram_w16_l512_id9_1_0_wenable;
  wire ram_w16_l512_id9_1_0_enable;
  wire [8-1:0] ram_w16_l512_id9_1_1_addr;
  wire [16-1:0] ram_w16_l512_id9_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id9_1_1_wdata;
  wire ram_w16_l512_id9_1_1_wenable;
  wire ram_w16_l512_id9_1_1_enable;
  assign ram_w16_l512_id9_1_0_wdata = 'hx;
  assign ram_w16_l512_id9_1_0_wenable = 0;

  ram_w16_l512_id9_1
  inst_ram_w16_l512_id9_1
  (
    .CLK(CLK),
    .ram_w16_l512_id9_1_0_addr(ram_w16_l512_id9_1_0_addr),
    .ram_w16_l512_id9_1_0_rdata(ram_w16_l512_id9_1_0_rdata),
    .ram_w16_l512_id9_1_0_wdata(ram_w16_l512_id9_1_0_wdata),
    .ram_w16_l512_id9_1_0_wenable(ram_w16_l512_id9_1_0_wenable),
    .ram_w16_l512_id9_1_0_enable(ram_w16_l512_id9_1_0_enable),
    .ram_w16_l512_id9_1_1_addr(ram_w16_l512_id9_1_1_addr),
    .ram_w16_l512_id9_1_1_rdata(ram_w16_l512_id9_1_1_rdata),
    .ram_w16_l512_id9_1_1_wdata(ram_w16_l512_id9_1_1_wdata),
    .ram_w16_l512_id9_1_1_wenable(ram_w16_l512_id9_1_1_wenable),
    .ram_w16_l512_id9_1_1_enable(ram_w16_l512_id9_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id10_0_0_addr;
  wire [16-1:0] ram_w16_l512_id10_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id10_0_0_wdata;
  wire ram_w16_l512_id10_0_0_wenable;
  wire ram_w16_l512_id10_0_0_enable;
  wire [8-1:0] ram_w16_l512_id10_0_1_addr;
  wire [16-1:0] ram_w16_l512_id10_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id10_0_1_wdata;
  wire ram_w16_l512_id10_0_1_wenable;
  wire ram_w16_l512_id10_0_1_enable;
  assign ram_w16_l512_id10_0_0_wdata = 'hx;
  assign ram_w16_l512_id10_0_0_wenable = 0;

  ram_w16_l512_id10_0
  inst_ram_w16_l512_id10_0
  (
    .CLK(CLK),
    .ram_w16_l512_id10_0_0_addr(ram_w16_l512_id10_0_0_addr),
    .ram_w16_l512_id10_0_0_rdata(ram_w16_l512_id10_0_0_rdata),
    .ram_w16_l512_id10_0_0_wdata(ram_w16_l512_id10_0_0_wdata),
    .ram_w16_l512_id10_0_0_wenable(ram_w16_l512_id10_0_0_wenable),
    .ram_w16_l512_id10_0_0_enable(ram_w16_l512_id10_0_0_enable),
    .ram_w16_l512_id10_0_1_addr(ram_w16_l512_id10_0_1_addr),
    .ram_w16_l512_id10_0_1_rdata(ram_w16_l512_id10_0_1_rdata),
    .ram_w16_l512_id10_0_1_wdata(ram_w16_l512_id10_0_1_wdata),
    .ram_w16_l512_id10_0_1_wenable(ram_w16_l512_id10_0_1_wenable),
    .ram_w16_l512_id10_0_1_enable(ram_w16_l512_id10_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id10_1_0_addr;
  wire [16-1:0] ram_w16_l512_id10_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id10_1_0_wdata;
  wire ram_w16_l512_id10_1_0_wenable;
  wire ram_w16_l512_id10_1_0_enable;
  wire [8-1:0] ram_w16_l512_id10_1_1_addr;
  wire [16-1:0] ram_w16_l512_id10_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id10_1_1_wdata;
  wire ram_w16_l512_id10_1_1_wenable;
  wire ram_w16_l512_id10_1_1_enable;
  assign ram_w16_l512_id10_1_0_wdata = 'hx;
  assign ram_w16_l512_id10_1_0_wenable = 0;

  ram_w16_l512_id10_1
  inst_ram_w16_l512_id10_1
  (
    .CLK(CLK),
    .ram_w16_l512_id10_1_0_addr(ram_w16_l512_id10_1_0_addr),
    .ram_w16_l512_id10_1_0_rdata(ram_w16_l512_id10_1_0_rdata),
    .ram_w16_l512_id10_1_0_wdata(ram_w16_l512_id10_1_0_wdata),
    .ram_w16_l512_id10_1_0_wenable(ram_w16_l512_id10_1_0_wenable),
    .ram_w16_l512_id10_1_0_enable(ram_w16_l512_id10_1_0_enable),
    .ram_w16_l512_id10_1_1_addr(ram_w16_l512_id10_1_1_addr),
    .ram_w16_l512_id10_1_1_rdata(ram_w16_l512_id10_1_1_rdata),
    .ram_w16_l512_id10_1_1_wdata(ram_w16_l512_id10_1_1_wdata),
    .ram_w16_l512_id10_1_1_wenable(ram_w16_l512_id10_1_1_wenable),
    .ram_w16_l512_id10_1_1_enable(ram_w16_l512_id10_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id11_0_0_addr;
  wire [16-1:0] ram_w16_l512_id11_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id11_0_0_wdata;
  wire ram_w16_l512_id11_0_0_wenable;
  wire ram_w16_l512_id11_0_0_enable;
  wire [8-1:0] ram_w16_l512_id11_0_1_addr;
  wire [16-1:0] ram_w16_l512_id11_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id11_0_1_wdata;
  wire ram_w16_l512_id11_0_1_wenable;
  wire ram_w16_l512_id11_0_1_enable;
  assign ram_w16_l512_id11_0_0_wdata = 'hx;
  assign ram_w16_l512_id11_0_0_wenable = 0;

  ram_w16_l512_id11_0
  inst_ram_w16_l512_id11_0
  (
    .CLK(CLK),
    .ram_w16_l512_id11_0_0_addr(ram_w16_l512_id11_0_0_addr),
    .ram_w16_l512_id11_0_0_rdata(ram_w16_l512_id11_0_0_rdata),
    .ram_w16_l512_id11_0_0_wdata(ram_w16_l512_id11_0_0_wdata),
    .ram_w16_l512_id11_0_0_wenable(ram_w16_l512_id11_0_0_wenable),
    .ram_w16_l512_id11_0_0_enable(ram_w16_l512_id11_0_0_enable),
    .ram_w16_l512_id11_0_1_addr(ram_w16_l512_id11_0_1_addr),
    .ram_w16_l512_id11_0_1_rdata(ram_w16_l512_id11_0_1_rdata),
    .ram_w16_l512_id11_0_1_wdata(ram_w16_l512_id11_0_1_wdata),
    .ram_w16_l512_id11_0_1_wenable(ram_w16_l512_id11_0_1_wenable),
    .ram_w16_l512_id11_0_1_enable(ram_w16_l512_id11_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id11_1_0_addr;
  wire [16-1:0] ram_w16_l512_id11_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id11_1_0_wdata;
  wire ram_w16_l512_id11_1_0_wenable;
  wire ram_w16_l512_id11_1_0_enable;
  wire [8-1:0] ram_w16_l512_id11_1_1_addr;
  wire [16-1:0] ram_w16_l512_id11_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id11_1_1_wdata;
  wire ram_w16_l512_id11_1_1_wenable;
  wire ram_w16_l512_id11_1_1_enable;
  assign ram_w16_l512_id11_1_0_wdata = 'hx;
  assign ram_w16_l512_id11_1_0_wenable = 0;

  ram_w16_l512_id11_1
  inst_ram_w16_l512_id11_1
  (
    .CLK(CLK),
    .ram_w16_l512_id11_1_0_addr(ram_w16_l512_id11_1_0_addr),
    .ram_w16_l512_id11_1_0_rdata(ram_w16_l512_id11_1_0_rdata),
    .ram_w16_l512_id11_1_0_wdata(ram_w16_l512_id11_1_0_wdata),
    .ram_w16_l512_id11_1_0_wenable(ram_w16_l512_id11_1_0_wenable),
    .ram_w16_l512_id11_1_0_enable(ram_w16_l512_id11_1_0_enable),
    .ram_w16_l512_id11_1_1_addr(ram_w16_l512_id11_1_1_addr),
    .ram_w16_l512_id11_1_1_rdata(ram_w16_l512_id11_1_1_rdata),
    .ram_w16_l512_id11_1_1_wdata(ram_w16_l512_id11_1_1_wdata),
    .ram_w16_l512_id11_1_1_wenable(ram_w16_l512_id11_1_1_wenable),
    .ram_w16_l512_id11_1_1_enable(ram_w16_l512_id11_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id12_0_0_addr;
  wire [16-1:0] ram_w16_l512_id12_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id12_0_0_wdata;
  wire ram_w16_l512_id12_0_0_wenable;
  wire ram_w16_l512_id12_0_0_enable;
  wire [8-1:0] ram_w16_l512_id12_0_1_addr;
  wire [16-1:0] ram_w16_l512_id12_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id12_0_1_wdata;
  wire ram_w16_l512_id12_0_1_wenable;
  wire ram_w16_l512_id12_0_1_enable;
  assign ram_w16_l512_id12_0_0_addr = 'hx;
  assign ram_w16_l512_id12_0_0_wdata = 'hx;
  assign ram_w16_l512_id12_0_0_wenable = 0;
  assign ram_w16_l512_id12_0_0_enable = 0;
  assign ram_w16_l512_id12_0_1_addr = 'hx;
  assign ram_w16_l512_id12_0_1_wdata = 'hx;
  assign ram_w16_l512_id12_0_1_wenable = 0;
  assign ram_w16_l512_id12_0_1_enable = 0;

  ram_w16_l512_id12_0
  inst_ram_w16_l512_id12_0
  (
    .CLK(CLK),
    .ram_w16_l512_id12_0_0_addr(ram_w16_l512_id12_0_0_addr),
    .ram_w16_l512_id12_0_0_rdata(ram_w16_l512_id12_0_0_rdata),
    .ram_w16_l512_id12_0_0_wdata(ram_w16_l512_id12_0_0_wdata),
    .ram_w16_l512_id12_0_0_wenable(ram_w16_l512_id12_0_0_wenable),
    .ram_w16_l512_id12_0_0_enable(ram_w16_l512_id12_0_0_enable),
    .ram_w16_l512_id12_0_1_addr(ram_w16_l512_id12_0_1_addr),
    .ram_w16_l512_id12_0_1_rdata(ram_w16_l512_id12_0_1_rdata),
    .ram_w16_l512_id12_0_1_wdata(ram_w16_l512_id12_0_1_wdata),
    .ram_w16_l512_id12_0_1_wenable(ram_w16_l512_id12_0_1_wenable),
    .ram_w16_l512_id12_0_1_enable(ram_w16_l512_id12_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id12_1_0_addr;
  wire [16-1:0] ram_w16_l512_id12_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id12_1_0_wdata;
  wire ram_w16_l512_id12_1_0_wenable;
  wire ram_w16_l512_id12_1_0_enable;
  wire [8-1:0] ram_w16_l512_id12_1_1_addr;
  wire [16-1:0] ram_w16_l512_id12_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id12_1_1_wdata;
  wire ram_w16_l512_id12_1_1_wenable;
  wire ram_w16_l512_id12_1_1_enable;
  assign ram_w16_l512_id12_1_0_addr = 'hx;
  assign ram_w16_l512_id12_1_0_wdata = 'hx;
  assign ram_w16_l512_id12_1_0_wenable = 0;
  assign ram_w16_l512_id12_1_0_enable = 0;
  assign ram_w16_l512_id12_1_1_addr = 'hx;
  assign ram_w16_l512_id12_1_1_wdata = 'hx;
  assign ram_w16_l512_id12_1_1_wenable = 0;
  assign ram_w16_l512_id12_1_1_enable = 0;

  ram_w16_l512_id12_1
  inst_ram_w16_l512_id12_1
  (
    .CLK(CLK),
    .ram_w16_l512_id12_1_0_addr(ram_w16_l512_id12_1_0_addr),
    .ram_w16_l512_id12_1_0_rdata(ram_w16_l512_id12_1_0_rdata),
    .ram_w16_l512_id12_1_0_wdata(ram_w16_l512_id12_1_0_wdata),
    .ram_w16_l512_id12_1_0_wenable(ram_w16_l512_id12_1_0_wenable),
    .ram_w16_l512_id12_1_0_enable(ram_w16_l512_id12_1_0_enable),
    .ram_w16_l512_id12_1_1_addr(ram_w16_l512_id12_1_1_addr),
    .ram_w16_l512_id12_1_1_rdata(ram_w16_l512_id12_1_1_rdata),
    .ram_w16_l512_id12_1_1_wdata(ram_w16_l512_id12_1_1_wdata),
    .ram_w16_l512_id12_1_1_wenable(ram_w16_l512_id12_1_1_wenable),
    .ram_w16_l512_id12_1_1_enable(ram_w16_l512_id12_1_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id0_0_addr;
  wire [32-1:0] ram_w32_l128_id0_0_rdata;
  wire [32-1:0] ram_w32_l128_id0_0_wdata;
  wire ram_w32_l128_id0_0_wenable;
  wire ram_w32_l128_id0_0_enable;
  wire [7-1:0] ram_w32_l128_id0_1_addr;
  wire [32-1:0] ram_w32_l128_id0_1_rdata;
  wire [32-1:0] ram_w32_l128_id0_1_wdata;
  wire ram_w32_l128_id0_1_wenable;
  wire ram_w32_l128_id0_1_enable;
  assign ram_w32_l128_id0_1_wdata = 'hx;
  assign ram_w32_l128_id0_1_wenable = 0;

  ram_w32_l128_id0
  inst_ram_w32_l128_id0
  (
    .CLK(CLK),
    .ram_w32_l128_id0_0_addr(ram_w32_l128_id0_0_addr),
    .ram_w32_l128_id0_0_rdata(ram_w32_l128_id0_0_rdata),
    .ram_w32_l128_id0_0_wdata(ram_w32_l128_id0_0_wdata),
    .ram_w32_l128_id0_0_wenable(ram_w32_l128_id0_0_wenable),
    .ram_w32_l128_id0_0_enable(ram_w32_l128_id0_0_enable),
    .ram_w32_l128_id0_1_addr(ram_w32_l128_id0_1_addr),
    .ram_w32_l128_id0_1_rdata(ram_w32_l128_id0_1_rdata),
    .ram_w32_l128_id0_1_wdata(ram_w32_l128_id0_1_wdata),
    .ram_w32_l128_id0_1_wenable(ram_w32_l128_id0_1_wenable),
    .ram_w32_l128_id0_1_enable(ram_w32_l128_id0_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id1_0_addr;
  wire [32-1:0] ram_w32_l128_id1_0_rdata;
  wire [32-1:0] ram_w32_l128_id1_0_wdata;
  wire ram_w32_l128_id1_0_wenable;
  wire ram_w32_l128_id1_0_enable;
  wire [7-1:0] ram_w32_l128_id1_1_addr;
  wire [32-1:0] ram_w32_l128_id1_1_rdata;
  wire [32-1:0] ram_w32_l128_id1_1_wdata;
  wire ram_w32_l128_id1_1_wenable;
  wire ram_w32_l128_id1_1_enable;
  assign ram_w32_l128_id1_0_wdata = 'hx;
  assign ram_w32_l128_id1_0_wenable = 0;

  ram_w32_l128_id1
  inst_ram_w32_l128_id1
  (
    .CLK(CLK),
    .ram_w32_l128_id1_0_addr(ram_w32_l128_id1_0_addr),
    .ram_w32_l128_id1_0_rdata(ram_w32_l128_id1_0_rdata),
    .ram_w32_l128_id1_0_wdata(ram_w32_l128_id1_0_wdata),
    .ram_w32_l128_id1_0_wenable(ram_w32_l128_id1_0_wenable),
    .ram_w32_l128_id1_0_enable(ram_w32_l128_id1_0_enable),
    .ram_w32_l128_id1_1_addr(ram_w32_l128_id1_1_addr),
    .ram_w32_l128_id1_1_rdata(ram_w32_l128_id1_1_rdata),
    .ram_w32_l128_id1_1_wdata(ram_w32_l128_id1_1_wdata),
    .ram_w32_l128_id1_1_wenable(ram_w32_l128_id1_1_wenable),
    .ram_w32_l128_id1_1_enable(ram_w32_l128_id1_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id2_0_addr;
  wire [32-1:0] ram_w32_l128_id2_0_rdata;
  wire [32-1:0] ram_w32_l128_id2_0_wdata;
  wire ram_w32_l128_id2_0_wenable;
  wire ram_w32_l128_id2_0_enable;
  wire [7-1:0] ram_w32_l128_id2_1_addr;
  wire [32-1:0] ram_w32_l128_id2_1_rdata;
  wire [32-1:0] ram_w32_l128_id2_1_wdata;
  wire ram_w32_l128_id2_1_wenable;
  wire ram_w32_l128_id2_1_enable;
  assign ram_w32_l128_id2_0_wdata = 'hx;
  assign ram_w32_l128_id2_0_wenable = 0;

  ram_w32_l128_id2
  inst_ram_w32_l128_id2
  (
    .CLK(CLK),
    .ram_w32_l128_id2_0_addr(ram_w32_l128_id2_0_addr),
    .ram_w32_l128_id2_0_rdata(ram_w32_l128_id2_0_rdata),
    .ram_w32_l128_id2_0_wdata(ram_w32_l128_id2_0_wdata),
    .ram_w32_l128_id2_0_wenable(ram_w32_l128_id2_0_wenable),
    .ram_w32_l128_id2_0_enable(ram_w32_l128_id2_0_enable),
    .ram_w32_l128_id2_1_addr(ram_w32_l128_id2_1_addr),
    .ram_w32_l128_id2_1_rdata(ram_w32_l128_id2_1_rdata),
    .ram_w32_l128_id2_1_wdata(ram_w32_l128_id2_1_wdata),
    .ram_w32_l128_id2_1_wenable(ram_w32_l128_id2_1_wenable),
    .ram_w32_l128_id2_1_enable(ram_w32_l128_id2_1_enable)
  );

  wire [6-1:0] cparam_conv2d_4_act_num_col;
  wire [6-1:0] cparam_conv2d_4_act_num_row;
  wire [9-1:0] cparam_conv2d_4_filter_num_och;
  wire [1-1:0] cparam_conv2d_4_bias_scala;
  wire [9-1:0] cparam_conv2d_4_bias_num;
  wire [1-1:0] cparam_conv2d_4_scale_scala;
  wire [9-1:0] cparam_conv2d_4_scale_num;
  wire [1-1:0] cparam_conv2d_4_vshamt_mul_scala;
  wire [1-1:0] cparam_conv2d_4_vshamt_mul_num;
  wire [1-1:0] cparam_conv2d_4_vshamt_sum_scala;
  wire [1-1:0] cparam_conv2d_4_vshamt_sum_num;
  wire [1-1:0] cparam_conv2d_4_vshamt_out_scala;
  wire [1-1:0] cparam_conv2d_4_vshamt_out_num;
  wire [1-1:0] cparam_conv2d_4_cshamt_mul_value;
  wire [1-1:0] cparam_conv2d_4_cshamt_sum_value;
  wire [1-1:0] cparam_conv2d_4_cshamt_out_value;
  wire [1-1:0] cparam_conv2d_4_act_func_index;
  wire [6-1:0] cparam_conv2d_4_out_num_col;
  wire [6-1:0] cparam_conv2d_4_out_num_row;
  wire [1-1:0] cparam_conv2d_4_pad_col_left;
  wire [1-1:0] cparam_conv2d_4_pad_row_top;
  wire [5-1:0] cparam_conv2d_4_max_col_count;
  wire [5-1:0] cparam_conv2d_4_max_row_count;
  wire [1-1:0] cparam_conv2d_4_max_bat_count;
  wire [8-1:0] cparam_conv2d_4_max_och_count;
  wire [4-1:0] cparam_conv2d_4_och_count_step;
  wire [1-1:0] cparam_conv2d_4_dma_flag_conds_0;
  wire [1-1:0] cparam_conv2d_4_dma_flag_conds_1;
  wire [1-1:0] cparam_conv2d_4_dma_flag_conds_2;
  wire signed [32-1:0] cparam_conv2d_4_act_offset_values_0;
  wire signed [32-1:0] cparam_conv2d_4_act_offset_values_1;
  wire signed [32-1:0] cparam_conv2d_4_act_offset_values_2;
  wire [12-1:0] cparam_conv2d_4_act_row_step;
  wire [16-1:0] cparam_conv2d_4_act_bat_step;
  wire [11-1:0] cparam_conv2d_4_act_read_size;
  wire [8-1:0] cparam_conv2d_4_act_read_block;
  wire [9-1:0] cparam_conv2d_4_act_read_step;
  wire [13-1:0] cparam_conv2d_4_filter_base_step;
  wire [12-1:0] cparam_conv2d_4_filter_read_size;
  wire [8-1:0] cparam_conv2d_4_filter_read_block;
  wire [9-1:0] cparam_conv2d_4_filter_read_step;
  wire [1-1:0] cparam_conv2d_4_out_offset_values_0;
  wire [10-1:0] cparam_conv2d_4_out_col_step;
  wire [13-1:0] cparam_conv2d_4_out_row_step;
  wire [18-1:0] cparam_conv2d_4_out_bat_step;
  wire [5-1:0] cparam_conv2d_4_out_och_step;
  wire [4-1:0] cparam_conv2d_4_out_write_size;
  wire [4-1:0] cparam_conv2d_4_out_write_size_res;
  wire [1-1:0] cparam_conv2d_4_out_write_block;
  wire [1-1:0] cparam_conv2d_4_keep_filter;
  wire [1-1:0] cparam_conv2d_4_keep_input;
  wire [1-1:0] cparam_conv2d_4_data_stationary;
  wire [4-1:0] cparam_conv2d_4_stream_num_ops;
  wire [4-1:0] cparam_conv2d_4_stream_num_ops_res;
  wire [4-1:0] cparam_conv2d_4_stream_num_ops_par;
  wire [4-1:0] cparam_conv2d_4_stream_num_ops_res_par;
  wire [8-1:0] cparam_conv2d_4_stream_reduce_size;
  wire [8-1:0] cparam_conv2d_4_stream_aligned_reduce_size;
  wire [1-1:0] cparam_conv2d_4_stream_omit_mask;
  wire [2-1:0] cparam_conv2d_4_col_select_initval;
  wire [1-1:0] cparam_conv2d_4_stride_col_par_col;
  wire [1-1:0] cparam_conv2d_4_stride_row_par_row;
  wire [1-1:0] cparam_conv2d_4_stride_col_mod_filter_num;
  wire [2-1:0] cparam_conv2d_4_filter_num_col_minus_stride_col_mod;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_0;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_1;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_2;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_3;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_4;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_5;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_6;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_7;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_8;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_9;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_10;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_11;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_12;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_13;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_14;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_15;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_16;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_17;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_18;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_19;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_20;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_21;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_22;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_23;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_24;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_25;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_26;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_small;
  wire [8-1:0] cparam_conv2d_4_inc_act_laddr_large;
  wire [9-1:0] cparam_conv2d_4_inc_out_laddr_col;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_small_offset;
  wire signed [9-1:0] cparam_conv2d_4_stream_act_local_large_offset;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_small_flags_1;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_small_flags_2;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_large_flags_1;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_large_flags_2;
  wire [1-1:0] cparam_conv2d_4_inc_sync_out;
  wire [1-1:0] cparam_conv2d_4_inc_sync_out_res;
  reg [2-1:0] conv2d_4_control_param_index;
  assign cparam_conv2d_4_act_num_col = (conv2d_4_control_param_index == 0)? 32'h20 : 
                                       (conv2d_4_control_param_index == 1)? 32'h10 : 32'h8;
  assign cparam_conv2d_4_act_num_row = (conv2d_4_control_param_index == 0)? 32'h20 : 
                                       (conv2d_4_control_param_index == 1)? 32'h10 : 32'h8;
  assign cparam_conv2d_4_filter_num_och = (conv2d_4_control_param_index == 0)? 32'h40 : 
                                          (conv2d_4_control_param_index == 1)? 32'h80 : 32'h100;
  assign cparam_conv2d_4_bias_scala = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                      (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_bias_num = (conv2d_4_control_param_index == 0)? 32'h40 : 
                                    (conv2d_4_control_param_index == 1)? 32'h80 : 32'h100;
  assign cparam_conv2d_4_scale_scala = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                       (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_scale_num = (conv2d_4_control_param_index == 0)? 32'h40 : 
                                     (conv2d_4_control_param_index == 1)? 32'h80 : 32'h100;
  assign cparam_conv2d_4_vshamt_mul_scala = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                            (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_vshamt_mul_num = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                          (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_vshamt_sum_scala = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                            (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_vshamt_sum_num = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                          (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_vshamt_out_scala = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                            (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_vshamt_out_num = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                          (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_cshamt_mul_value = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                            (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_cshamt_sum_value = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                            (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_cshamt_out_value = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                            (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_act_func_index = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                          (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_out_num_col = (conv2d_4_control_param_index == 0)? 32'h20 : 
                                       (conv2d_4_control_param_index == 1)? 32'h10 : 32'h8;
  assign cparam_conv2d_4_out_num_row = (conv2d_4_control_param_index == 0)? 32'h20 : 
                                       (conv2d_4_control_param_index == 1)? 32'h10 : 32'h8;
  assign cparam_conv2d_4_pad_col_left = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                        (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_pad_row_top = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                       (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_max_col_count = (conv2d_4_control_param_index == 0)? 32'h1f : 
                                         (conv2d_4_control_param_index == 1)? 32'hf : 32'h7;
  assign cparam_conv2d_4_max_row_count = (conv2d_4_control_param_index == 0)? 32'h1f : 
                                         (conv2d_4_control_param_index == 1)? 32'hf : 32'h7;
  assign cparam_conv2d_4_max_bat_count = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                         (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_max_och_count = (conv2d_4_control_param_index == 0)? 32'h38 : 
                                         (conv2d_4_control_param_index == 1)? 32'h7c : 32'hfe;
  assign cparam_conv2d_4_och_count_step = (conv2d_4_control_param_index == 0)? 32'h8 : 
                                          (conv2d_4_control_param_index == 1)? 32'h4 : 32'h2;
  assign cparam_conv2d_4_dma_flag_conds_0 = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                            (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_dma_flag_conds_1 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                            (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_dma_flag_conds_2 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                            (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_act_offset_values_0 = (conv2d_4_control_param_index == 0)? -32'sh100 : 
                                               (conv2d_4_control_param_index == 1)? -32'sh800 : -32'sh800;
  assign cparam_conv2d_4_act_offset_values_1 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                               (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_act_offset_values_2 = (conv2d_4_control_param_index == 0)? 32'h100 : 
                                               (conv2d_4_control_param_index == 1)? 32'h800 : 32'h800;
  assign cparam_conv2d_4_act_row_step = (conv2d_4_control_param_index == 0)? 32'h100 : 
                                        (conv2d_4_control_param_index == 1)? 32'h800 : 32'h800;
  assign cparam_conv2d_4_act_bat_step = (conv2d_4_control_param_index == 0)? 32'h2000 : 
                                        (conv2d_4_control_param_index == 1)? 32'h8000 : 32'h4000;
  assign cparam_conv2d_4_act_read_size = (conv2d_4_control_param_index == 0)? 32'h80 : 
                                         (conv2d_4_control_param_index == 1)? 32'h400 : 32'h400;
  assign cparam_conv2d_4_act_read_block = (conv2d_4_control_param_index == 0)? 32'h4 : 
                                          (conv2d_4_control_param_index == 1)? 32'h40 : 32'h80;
  assign cparam_conv2d_4_act_read_step = (conv2d_4_control_param_index == 0)? 32'h2c : 
                                         (conv2d_4_control_param_index == 1)? 32'h180 : 32'h180;
  assign cparam_conv2d_4_filter_base_step = (conv2d_4_control_param_index == 0)? 32'h240 : 
                                            (conv2d_4_control_param_index == 1)? 32'h1200 : 32'h1200;
  assign cparam_conv2d_4_filter_read_size = (conv2d_4_control_param_index == 0)? 32'h120 : 
                                            (conv2d_4_control_param_index == 1)? 32'h900 : 32'h900;
  assign cparam_conv2d_4_filter_read_block = (conv2d_4_control_param_index == 0)? 32'h4 : 
                                             (conv2d_4_control_param_index == 1)? 32'h40 : 32'h80;
  assign cparam_conv2d_4_filter_read_step = (conv2d_4_control_param_index == 0)? 32'h20 : 
                                            (conv2d_4_control_param_index == 1)? 32'h100 : 32'h100;
  assign cparam_conv2d_4_out_offset_values_0 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                               (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_out_col_step = (conv2d_4_control_param_index == 0)? 32'h80 : 
                                        (conv2d_4_control_param_index == 1)? 32'h100 : 32'h200;
  assign cparam_conv2d_4_out_row_step = (conv2d_4_control_param_index == 0)? 32'h1000 : 
                                        (conv2d_4_control_param_index == 1)? 32'h1000 : 32'h1000;
  assign cparam_conv2d_4_out_bat_step = (conv2d_4_control_param_index == 0)? 32'h20000 : 
                                        (conv2d_4_control_param_index == 1)? 32'h10000 : 32'h8000;
  assign cparam_conv2d_4_out_och_step = (conv2d_4_control_param_index == 0)? 32'h10 : 
                                        (conv2d_4_control_param_index == 1)? 32'h8 : 32'h4;
  assign cparam_conv2d_4_out_write_size = (conv2d_4_control_param_index == 0)? 32'h8 : 
                                          (conv2d_4_control_param_index == 1)? 32'h4 : 32'h2;
  assign cparam_conv2d_4_out_write_size_res = (conv2d_4_control_param_index == 0)? 32'h8 : 
                                              (conv2d_4_control_param_index == 1)? 32'h4 : 32'h2;
  assign cparam_conv2d_4_out_write_block = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                           (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_keep_filter = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                       (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_keep_input = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                      (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_data_stationary = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                           (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_stream_num_ops = (conv2d_4_control_param_index == 0)? 32'h8 : 
                                          (conv2d_4_control_param_index == 1)? 32'h4 : 32'h2;
  assign cparam_conv2d_4_stream_num_ops_res = (conv2d_4_control_param_index == 0)? 32'h8 : 
                                              (conv2d_4_control_param_index == 1)? 32'h4 : 32'h2;
  assign cparam_conv2d_4_stream_num_ops_par = (conv2d_4_control_param_index == 0)? 32'h8 : 
                                              (conv2d_4_control_param_index == 1)? 32'h4 : 32'h2;
  assign cparam_conv2d_4_stream_num_ops_res_par = (conv2d_4_control_param_index == 0)? 32'h8 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h4 : 32'h2;
  assign cparam_conv2d_4_stream_reduce_size = (conv2d_4_control_param_index == 0)? 32'h3 : 
                                              (conv2d_4_control_param_index == 1)? 32'h40 : 32'h80;
  assign cparam_conv2d_4_stream_aligned_reduce_size = (conv2d_4_control_param_index == 0)? 32'h4 : 
                                                      (conv2d_4_control_param_index == 1)? 32'h40 : 32'h80;
  assign cparam_conv2d_4_stream_omit_mask = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                            (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_col_select_initval = (conv2d_4_control_param_index == 0)? 32'h2 : 
                                              (conv2d_4_control_param_index == 1)? 32'h2 : 32'h2;
  assign cparam_conv2d_4_stride_col_par_col = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                              (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_stride_row_par_row = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                              (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_stride_col_mod_filter_num = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                                     (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_filter_num_col_minus_stride_col_mod = (conv2d_4_control_param_index == 0)? 32'h2 : 
                                                               (conv2d_4_control_param_index == 1)? 32'h2 : 32'h2;
  assign cparam_conv2d_4_inc_act_laddr_conds_0 = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                                 (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_1 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                 (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_2 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                 (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_3 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                 (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_4 = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                                 (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_5 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                 (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_6 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                 (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_7 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                 (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_8 = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                                 (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_9 = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                                 (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_10 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_11 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_12 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_13 = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_14 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_15 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_16 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_17 = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_18 = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_19 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_20 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_21 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_22 = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_23 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_24 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_25 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_26 = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                                  (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_small = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                               (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_large = (conv2d_4_control_param_index == 0)? 32'h4 : 
                                               (conv2d_4_control_param_index == 1)? 32'h40 : 32'h80;
  assign cparam_conv2d_4_inc_out_laddr_col = (conv2d_4_control_param_index == 0)? 32'h40 : 
                                             (conv2d_4_control_param_index == 1)? 32'h80 : 32'h100;
  assign cparam_conv2d_4_stream_act_local_small_offset = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                         (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_stream_act_local_large_offset = (conv2d_4_control_param_index == 0)? -32'sh4 : 
                                                         (conv2d_4_control_param_index == 1)? -32'sh40 : -32'sh80;
  assign cparam_conv2d_4_stream_act_local_small_flags_0 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                          (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_stream_act_local_small_flags_1 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                          (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_stream_act_local_small_flags_2 = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                                          (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_stream_act_local_large_flags_0 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                          (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_stream_act_local_large_flags_1 = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                                          (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_stream_act_local_large_flags_2 = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                                          (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_sync_out = (conv2d_4_control_param_index == 0)? 32'h1 : 
                                        (conv2d_4_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_sync_out_res = (conv2d_4_control_param_index == 0)? 32'h0 : 
                                            (conv2d_4_control_param_index == 1)? 32'h0 : 32'h0;
  wire [6-1:0] cparam_max_pool_serial_6_act_num_col;
  wire [6-1:0] cparam_max_pool_serial_6_act_num_row;
  wire [2-1:0] cparam_max_pool_serial_6_stride_col;
  wire [2-1:0] cparam_max_pool_serial_6_stride_row;
  wire [5-1:0] cparam_max_pool_serial_6_out_num_col;
  wire [5-1:0] cparam_max_pool_serial_6_out_num_row;
  wire [1-1:0] cparam_max_pool_serial_6_pad_col_left;
  wire [1-1:0] cparam_max_pool_serial_6_pad_row_top;
  wire [5-1:0] cparam_max_pool_serial_6_max_col_count;
  wire [5-1:0] cparam_max_pool_serial_6_max_row_count;
  wire [1-1:0] cparam_max_pool_serial_6_max_bat_count;
  wire signed [32-1:0] cparam_max_pool_serial_6_act_offset_values_0;
  wire signed [32-1:0] cparam_max_pool_serial_6_act_offset_values_1;
  wire [14-1:0] cparam_max_pool_serial_6_act_row_step;
  wire [18-1:0] cparam_max_pool_serial_6_act_bat_step;
  wire [11-1:0] cparam_max_pool_serial_6_act_read_size;
  wire [8-1:0] cparam_max_pool_serial_6_act_read_block;
  wire [12-1:0] cparam_max_pool_serial_6_out_row_step;
  wire [16-1:0] cparam_max_pool_serial_6_out_bat_step;
  wire [10-1:0] cparam_max_pool_serial_6_out_write_size;
  wire [8-1:0] cparam_max_pool_serial_6_stream_size;
  wire [1-1:0] cparam_max_pool_serial_6_col_select_initval;
  wire [1-1:0] cparam_max_pool_serial_6_stride_col_mod_ksize;
  wire [2-1:0] cparam_max_pool_serial_6_ksize_col_minus_stride_col_mod;
  wire [1-1:0] cparam_max_pool_serial_6_local_pad_offset;
  wire [9-1:0] cparam_max_pool_serial_6_inc_act_laddr;
  wire [8-1:0] cparam_max_pool_serial_6_inc_out_laddr;
  reg [2-1:0] max_pool_serial_6_control_param_index;
  assign cparam_max_pool_serial_6_act_num_col = (max_pool_serial_6_control_param_index == 0)? 32'h20 : 
                                                (max_pool_serial_6_control_param_index == 1)? 32'h10 : 32'h8;
  assign cparam_max_pool_serial_6_act_num_row = (max_pool_serial_6_control_param_index == 0)? 32'h20 : 
                                                (max_pool_serial_6_control_param_index == 1)? 32'h10 : 32'h8;
  assign cparam_max_pool_serial_6_stride_col = (max_pool_serial_6_control_param_index == 0)? 32'h2 : 
                                               (max_pool_serial_6_control_param_index == 1)? 32'h2 : 32'h2;
  assign cparam_max_pool_serial_6_stride_row = (max_pool_serial_6_control_param_index == 0)? 32'h2 : 
                                               (max_pool_serial_6_control_param_index == 1)? 32'h2 : 32'h2;
  assign cparam_max_pool_serial_6_out_num_col = (max_pool_serial_6_control_param_index == 0)? 32'h10 : 
                                                (max_pool_serial_6_control_param_index == 1)? 32'h8 : 32'h4;
  assign cparam_max_pool_serial_6_out_num_row = (max_pool_serial_6_control_param_index == 0)? 32'h10 : 
                                                (max_pool_serial_6_control_param_index == 1)? 32'h8 : 32'h4;
  assign cparam_max_pool_serial_6_pad_col_left = (max_pool_serial_6_control_param_index == 0)? 32'h0 : 
                                                 (max_pool_serial_6_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_6_pad_row_top = (max_pool_serial_6_control_param_index == 0)? 32'h0 : 
                                                (max_pool_serial_6_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_6_max_col_count = (max_pool_serial_6_control_param_index == 0)? 32'h1d : 
                                                  (max_pool_serial_6_control_param_index == 1)? 32'hd : 32'h5;
  assign cparam_max_pool_serial_6_max_row_count = (max_pool_serial_6_control_param_index == 0)? 32'h1d : 
                                                  (max_pool_serial_6_control_param_index == 1)? 32'hd : 32'h5;
  assign cparam_max_pool_serial_6_max_bat_count = (max_pool_serial_6_control_param_index == 0)? 32'h0 : 
                                                  (max_pool_serial_6_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_6_act_offset_values_0 = (max_pool_serial_6_control_param_index == 0)? 32'h0 : 
                                                        (max_pool_serial_6_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_6_act_offset_values_1 = (max_pool_serial_6_control_param_index == 0)? 32'h1000 : 
                                                        (max_pool_serial_6_control_param_index == 1)? 32'h1000 : 32'h1000;
  assign cparam_max_pool_serial_6_act_row_step = (max_pool_serial_6_control_param_index == 0)? 32'h2000 : 
                                                 (max_pool_serial_6_control_param_index == 1)? 32'h2000 : 32'h2000;
  assign cparam_max_pool_serial_6_act_bat_step = (max_pool_serial_6_control_param_index == 0)? 32'h20000 : 
                                                 (max_pool_serial_6_control_param_index == 1)? 32'h10000 : 32'h8000;
  assign cparam_max_pool_serial_6_act_read_size = (max_pool_serial_6_control_param_index == 0)? 32'h400 : 
                                                  (max_pool_serial_6_control_param_index == 1)? 32'h400 : 32'h400;
  assign cparam_max_pool_serial_6_act_read_block = (max_pool_serial_6_control_param_index == 0)? 32'h20 : 
                                                   (max_pool_serial_6_control_param_index == 1)? 32'h40 : 32'h80;
  assign cparam_max_pool_serial_6_out_row_step = (max_pool_serial_6_control_param_index == 0)? 32'h800 : 
                                                 (max_pool_serial_6_control_param_index == 1)? 32'h800 : 32'h800;
  assign cparam_max_pool_serial_6_out_bat_step = (max_pool_serial_6_control_param_index == 0)? 32'h8000 : 
                                                 (max_pool_serial_6_control_param_index == 1)? 32'h4000 : 32'h2000;
  assign cparam_max_pool_serial_6_out_write_size = (max_pool_serial_6_control_param_index == 0)? 32'h200 : 
                                                   (max_pool_serial_6_control_param_index == 1)? 32'h200 : 32'h200;
  assign cparam_max_pool_serial_6_stream_size = (max_pool_serial_6_control_param_index == 0)? 32'h20 : 
                                                (max_pool_serial_6_control_param_index == 1)? 32'h40 : 32'h80;
  assign cparam_max_pool_serial_6_col_select_initval = (max_pool_serial_6_control_param_index == 0)? 32'h0 : 
                                                       (max_pool_serial_6_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_6_stride_col_mod_ksize = (max_pool_serial_6_control_param_index == 0)? 32'h0 : 
                                                         (max_pool_serial_6_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_6_ksize_col_minus_stride_col_mod = (max_pool_serial_6_control_param_index == 0)? 32'h2 : 
                                                                   (max_pool_serial_6_control_param_index == 1)? 32'h2 : 32'h2;
  assign cparam_max_pool_serial_6_local_pad_offset = (max_pool_serial_6_control_param_index == 0)? 32'h0 : 
                                                     (max_pool_serial_6_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_6_inc_act_laddr = (max_pool_serial_6_control_param_index == 0)? 32'h40 : 
                                                  (max_pool_serial_6_control_param_index == 1)? 32'h80 : 32'h100;
  assign cparam_max_pool_serial_6_inc_out_laddr = (max_pool_serial_6_control_param_index == 0)? 32'h20 : 
                                                  (max_pool_serial_6_control_param_index == 1)? 32'h40 : 32'h80;
  wire [1-1:0] cparam_matmul_23_act_num_col;
  wire [1-1:0] cparam_matmul_23_act_num_row;
  wire [11-1:0] cparam_matmul_23_filter_num_och;
  wire [1-1:0] cparam_matmul_23_bias_scala;
  wire [11-1:0] cparam_matmul_23_bias_num;
  wire [1-1:0] cparam_matmul_23_scale_scala;
  wire [11-1:0] cparam_matmul_23_scale_num;
  wire [1-1:0] cparam_matmul_23_vshamt_mul_scala;
  wire [1-1:0] cparam_matmul_23_vshamt_mul_num;
  wire [1-1:0] cparam_matmul_23_vshamt_sum_scala;
  wire [1-1:0] cparam_matmul_23_vshamt_sum_num;
  wire [1-1:0] cparam_matmul_23_vshamt_out_scala;
  wire [1-1:0] cparam_matmul_23_vshamt_out_num;
  wire [1-1:0] cparam_matmul_23_cshamt_mul_value;
  wire [1-1:0] cparam_matmul_23_cshamt_sum_value;
  wire [1-1:0] cparam_matmul_23_cshamt_out_value;
  wire [1-1:0] cparam_matmul_23_act_func_index;
  wire [1-1:0] cparam_matmul_23_out_num_col;
  wire [1-1:0] cparam_matmul_23_out_num_row;
  wire [1-1:0] cparam_matmul_23_pad_col_left;
  wire [1-1:0] cparam_matmul_23_pad_row_top;
  wire [1-1:0] cparam_matmul_23_max_col_count;
  wire [1-1:0] cparam_matmul_23_max_row_count;
  wire [1-1:0] cparam_matmul_23_max_bat_count;
  wire [10-1:0] cparam_matmul_23_max_och_count;
  wire [4-1:0] cparam_matmul_23_och_count_step;
  wire [1-1:0] cparam_matmul_23_dma_flag_conds_0;
  wire signed [32-1:0] cparam_matmul_23_act_offset_values_0;
  wire [14-1:0] cparam_matmul_23_act_row_step;
  wire [14-1:0] cparam_matmul_23_act_bat_step;
  wire [13-1:0] cparam_matmul_23_act_read_size;
  wire [13-1:0] cparam_matmul_23_act_read_block;
  wire [13-1:0] cparam_matmul_23_act_read_step;
  wire [15-1:0] cparam_matmul_23_filter_base_step;
  wire [14-1:0] cparam_matmul_23_filter_read_size;
  wire [13-1:0] cparam_matmul_23_filter_read_block;
  wire [14-1:0] cparam_matmul_23_filter_read_step;
  wire [1-1:0] cparam_matmul_23_out_offset_values_0;
  wire [12-1:0] cparam_matmul_23_out_col_step;
  wire [12-1:0] cparam_matmul_23_out_row_step;
  wire [12-1:0] cparam_matmul_23_out_bat_step;
  wire [5-1:0] cparam_matmul_23_out_och_step;
  wire [4-1:0] cparam_matmul_23_out_write_size;
  wire [4-1:0] cparam_matmul_23_out_write_size_res;
  wire [1-1:0] cparam_matmul_23_out_write_block;
  wire [1-1:0] cparam_matmul_23_keep_filter;
  wire [1-1:0] cparam_matmul_23_keep_input;
  wire [1-1:0] cparam_matmul_23_data_stationary;
  wire [4-1:0] cparam_matmul_23_stream_num_ops;
  wire [4-1:0] cparam_matmul_23_stream_num_ops_res;
  wire [4-1:0] cparam_matmul_23_stream_num_ops_par;
  wire [4-1:0] cparam_matmul_23_stream_num_ops_res_par;
  wire [13-1:0] cparam_matmul_23_stream_reduce_size;
  wire [13-1:0] cparam_matmul_23_stream_aligned_reduce_size;
  wire [1-1:0] cparam_matmul_23_stream_omit_mask;
  wire [1-1:0] cparam_matmul_23_col_select_initval;
  wire [1-1:0] cparam_matmul_23_stride_col_par_col;
  wire [1-1:0] cparam_matmul_23_stride_row_par_row;
  wire [1-1:0] cparam_matmul_23_stride_col_mod_filter_num;
  wire [1-1:0] cparam_matmul_23_filter_num_col_minus_stride_col_mod;
  wire [1-1:0] cparam_matmul_23_inc_act_laddr_conds_0;
  wire [13-1:0] cparam_matmul_23_inc_act_laddr_small;
  wire [13-1:0] cparam_matmul_23_inc_act_laddr_large;
  wire [11-1:0] cparam_matmul_23_inc_out_laddr_col;
  wire [1-1:0] cparam_matmul_23_stream_act_local_small_offset;
  wire [1-1:0] cparam_matmul_23_stream_act_local_large_offset;
  wire [1-1:0] cparam_matmul_23_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_matmul_23_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_matmul_23_inc_sync_out;
  wire [1-1:0] cparam_matmul_23_inc_sync_out_res;
  reg [1-1:0] matmul_23_control_param_index;
  assign cparam_matmul_23_act_num_col = (matmul_23_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_23_act_num_row = (matmul_23_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_23_filter_num_och = (matmul_23_control_param_index == 0)? 32'h400 : 32'h200;
  assign cparam_matmul_23_bias_scala = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_bias_num = (matmul_23_control_param_index == 0)? 32'h400 : 32'h200;
  assign cparam_matmul_23_scale_scala = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_scale_num = (matmul_23_control_param_index == 0)? 32'h400 : 32'h200;
  assign cparam_matmul_23_vshamt_mul_scala = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_vshamt_mul_num = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_vshamt_sum_scala = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_vshamt_sum_num = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_vshamt_out_scala = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_vshamt_out_num = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_cshamt_mul_value = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_cshamt_sum_value = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_cshamt_out_value = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_act_func_index = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_out_num_col = (matmul_23_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_23_out_num_row = (matmul_23_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_23_pad_col_left = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_pad_row_top = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_max_col_count = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_max_row_count = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_max_bat_count = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_max_och_count = (matmul_23_control_param_index == 0)? 32'h3fe : 32'h1f8;
  assign cparam_matmul_23_och_count_step = (matmul_23_control_param_index == 0)? 32'h2 : 32'h8;
  assign cparam_matmul_23_dma_flag_conds_0 = (matmul_23_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_23_act_offset_values_0 = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_act_row_step = (matmul_23_control_param_index == 0)? 32'h2000 : 32'h800;
  assign cparam_matmul_23_act_bat_step = (matmul_23_control_param_index == 0)? 32'h2000 : 32'h800;
  assign cparam_matmul_23_act_read_size = (matmul_23_control_param_index == 0)? 32'h1000 : 32'h400;
  assign cparam_matmul_23_act_read_block = (matmul_23_control_param_index == 0)? 32'h1000 : 32'h400;
  assign cparam_matmul_23_act_read_step = (matmul_23_control_param_index == 0)? 32'h1000 : 32'h400;
  assign cparam_matmul_23_filter_base_step = (matmul_23_control_param_index == 0)? 32'h4000 : 32'h4000;
  assign cparam_matmul_23_filter_read_size = (matmul_23_control_param_index == 0)? 32'h2000 : 32'h2000;
  assign cparam_matmul_23_filter_read_block = (matmul_23_control_param_index == 0)? 32'h1000 : 32'h400;
  assign cparam_matmul_23_filter_read_step = (matmul_23_control_param_index == 0)? 32'h2000 : 32'h2000;
  assign cparam_matmul_23_out_offset_values_0 = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_out_col_step = (matmul_23_control_param_index == 0)? 32'h800 : 32'h400;
  assign cparam_matmul_23_out_row_step = (matmul_23_control_param_index == 0)? 32'h800 : 32'h400;
  assign cparam_matmul_23_out_bat_step = (matmul_23_control_param_index == 0)? 32'h800 : 32'h400;
  assign cparam_matmul_23_out_och_step = (matmul_23_control_param_index == 0)? 32'h4 : 32'h10;
  assign cparam_matmul_23_out_write_size = (matmul_23_control_param_index == 0)? 32'h2 : 32'h8;
  assign cparam_matmul_23_out_write_size_res = (matmul_23_control_param_index == 0)? 32'h2 : 32'h8;
  assign cparam_matmul_23_out_write_block = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_keep_filter = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_keep_input = (matmul_23_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_23_data_stationary = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_stream_num_ops = (matmul_23_control_param_index == 0)? 32'h2 : 32'h8;
  assign cparam_matmul_23_stream_num_ops_res = (matmul_23_control_param_index == 0)? 32'h2 : 32'h8;
  assign cparam_matmul_23_stream_num_ops_par = (matmul_23_control_param_index == 0)? 32'h2 : 32'h8;
  assign cparam_matmul_23_stream_num_ops_res_par = (matmul_23_control_param_index == 0)? 32'h2 : 32'h8;
  assign cparam_matmul_23_stream_reduce_size = (matmul_23_control_param_index == 0)? 32'h1000 : 32'h400;
  assign cparam_matmul_23_stream_aligned_reduce_size = (matmul_23_control_param_index == 0)? 32'h1000 : 32'h400;
  assign cparam_matmul_23_stream_omit_mask = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_col_select_initval = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_stride_col_par_col = (matmul_23_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_23_stride_row_par_row = (matmul_23_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_23_stride_col_mod_filter_num = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_filter_num_col_minus_stride_col_mod = (matmul_23_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_23_inc_act_laddr_conds_0 = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_inc_act_laddr_small = (matmul_23_control_param_index == 0)? 32'h1000 : 32'h400;
  assign cparam_matmul_23_inc_act_laddr_large = (matmul_23_control_param_index == 0)? 32'h1000 : 32'h400;
  assign cparam_matmul_23_inc_out_laddr_col = (matmul_23_control_param_index == 0)? 32'h400 : 32'h200;
  assign cparam_matmul_23_stream_act_local_small_offset = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_stream_act_local_large_offset = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_stream_act_local_small_flags_0 = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_stream_act_local_large_flags_0 = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_23_inc_sync_out = (matmul_23_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_23_inc_sync_out_res = (matmul_23_control_param_index == 0)? 32'h0 : 32'h0;
  wire [1-1:0] cparam_matmul_33_act_num_col;
  wire [1-1:0] cparam_matmul_33_act_num_row;
  wire [4-1:0] cparam_matmul_33_filter_num_och;
  wire [1-1:0] cparam_matmul_33_bias_scala;
  wire [3-1:0] cparam_matmul_33_bias_num;
  wire [1-1:0] cparam_matmul_33_scale_scala;
  wire [3-1:0] cparam_matmul_33_scale_num;
  wire [1-1:0] cparam_matmul_33_vshamt_mul_scala;
  wire [1-1:0] cparam_matmul_33_vshamt_mul_num;
  wire [1-1:0] cparam_matmul_33_vshamt_sum_scala;
  wire [1-1:0] cparam_matmul_33_vshamt_sum_num;
  wire [1-1:0] cparam_matmul_33_vshamt_out_scala;
  wire [1-1:0] cparam_matmul_33_vshamt_out_num;
  wire [1-1:0] cparam_matmul_33_cshamt_mul_value;
  wire [1-1:0] cparam_matmul_33_cshamt_sum_value;
  wire [5-1:0] cparam_matmul_33_cshamt_out_value;
  wire [1-1:0] cparam_matmul_33_act_func_index;
  wire [1-1:0] cparam_matmul_33_out_num_col;
  wire [1-1:0] cparam_matmul_33_out_num_row;
  wire [1-1:0] cparam_matmul_33_pad_col_left;
  wire [1-1:0] cparam_matmul_33_pad_row_top;
  wire [1-1:0] cparam_matmul_33_max_col_count;
  wire [1-1:0] cparam_matmul_33_max_row_count;
  wire [1-1:0] cparam_matmul_33_max_bat_count;
  wire [3-1:0] cparam_matmul_33_max_och_count;
  wire [1-1:0] cparam_matmul_33_och_count_step;
  wire [1-1:0] cparam_matmul_33_dma_flag_conds_0;
  wire signed [32-1:0] cparam_matmul_33_act_offset_values_0;
  wire [11-1:0] cparam_matmul_33_act_row_step;
  wire [11-1:0] cparam_matmul_33_act_bat_step;
  wire [9-1:0] cparam_matmul_33_act_read_size;
  wire [9-1:0] cparam_matmul_33_act_read_block;
  wire [9-1:0] cparam_matmul_33_act_read_step;
  wire [12-1:0] cparam_matmul_33_filter_base_step;
  wire [10-1:0] cparam_matmul_33_filter_read_size;
  wire [9-1:0] cparam_matmul_33_filter_read_block;
  wire [9-1:0] cparam_matmul_33_filter_read_step;
  wire [1-1:0] cparam_matmul_33_out_offset_values_0;
  wire [5-1:0] cparam_matmul_33_out_col_step;
  wire [5-1:0] cparam_matmul_33_out_row_step;
  wire [5-1:0] cparam_matmul_33_out_bat_step;
  wire [3-1:0] cparam_matmul_33_out_och_step;
  wire [1-1:0] cparam_matmul_33_out_write_size;
  wire [1-1:0] cparam_matmul_33_out_write_size_res;
  wire [1-1:0] cparam_matmul_33_out_write_block;
  wire [1-1:0] cparam_matmul_33_keep_filter;
  wire [1-1:0] cparam_matmul_33_keep_input;
  wire [1-1:0] cparam_matmul_33_data_stationary;
  wire [1-1:0] cparam_matmul_33_stream_num_ops;
  wire [1-1:0] cparam_matmul_33_stream_num_ops_res;
  wire [1-1:0] cparam_matmul_33_stream_num_ops_par;
  wire [1-1:0] cparam_matmul_33_stream_num_ops_res_par;
  wire [9-1:0] cparam_matmul_33_stream_reduce_size;
  wire [9-1:0] cparam_matmul_33_stream_aligned_reduce_size;
  wire [1-1:0] cparam_matmul_33_stream_omit_mask;
  wire [1-1:0] cparam_matmul_33_col_select_initval;
  wire [1-1:0] cparam_matmul_33_stride_col_par_col;
  wire [1-1:0] cparam_matmul_33_stride_row_par_row;
  wire [1-1:0] cparam_matmul_33_stride_col_mod_filter_num;
  wire [1-1:0] cparam_matmul_33_filter_num_col_minus_stride_col_mod;
  wire [1-1:0] cparam_matmul_33_inc_act_laddr_conds_0;
  wire [9-1:0] cparam_matmul_33_inc_act_laddr_small;
  wire [9-1:0] cparam_matmul_33_inc_act_laddr_large;
  wire [3-1:0] cparam_matmul_33_inc_out_laddr_col;
  wire [1-1:0] cparam_matmul_33_stream_act_local_small_offset;
  wire [1-1:0] cparam_matmul_33_stream_act_local_large_offset;
  wire [1-1:0] cparam_matmul_33_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_matmul_33_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_matmul_33_inc_sync_out;
  wire [1-1:0] cparam_matmul_33_inc_sync_out_res;
  assign cparam_matmul_33_act_num_col = 1;
  assign cparam_matmul_33_act_num_row = 1;
  assign cparam_matmul_33_filter_num_och = 10;
  assign cparam_matmul_33_bias_scala = 0;
  assign cparam_matmul_33_bias_num = 5;
  assign cparam_matmul_33_scale_scala = 0;
  assign cparam_matmul_33_scale_num = 5;
  assign cparam_matmul_33_vshamt_mul_scala = 0;
  assign cparam_matmul_33_vshamt_mul_num = 0;
  assign cparam_matmul_33_vshamt_sum_scala = 0;
  assign cparam_matmul_33_vshamt_sum_num = 0;
  assign cparam_matmul_33_vshamt_out_scala = 0;
  assign cparam_matmul_33_vshamt_out_num = 0;
  assign cparam_matmul_33_cshamt_mul_value = 0;
  assign cparam_matmul_33_cshamt_sum_value = 0;
  assign cparam_matmul_33_cshamt_out_value = 17;
  assign cparam_matmul_33_act_func_index = 0;
  assign cparam_matmul_33_out_num_col = 1;
  assign cparam_matmul_33_out_num_row = 1;
  assign cparam_matmul_33_pad_col_left = 0;
  assign cparam_matmul_33_pad_row_top = 0;
  assign cparam_matmul_33_max_col_count = 0;
  assign cparam_matmul_33_max_row_count = 0;
  assign cparam_matmul_33_max_bat_count = 0;
  assign cparam_matmul_33_max_och_count = 4;
  assign cparam_matmul_33_och_count_step = 1;
  assign cparam_matmul_33_dma_flag_conds_0 = 1;
  assign cparam_matmul_33_act_offset_values_0 = 0;
  assign cparam_matmul_33_act_row_step = 1024;
  assign cparam_matmul_33_act_bat_step = 1024;
  assign cparam_matmul_33_act_read_size = 256;
  assign cparam_matmul_33_act_read_block = 256;
  assign cparam_matmul_33_act_read_step = 256;
  assign cparam_matmul_33_filter_base_step = 2048;
  assign cparam_matmul_33_filter_read_size = 512;
  assign cparam_matmul_33_filter_read_block = 256;
  assign cparam_matmul_33_filter_read_step = 256;
  assign cparam_matmul_33_out_offset_values_0 = 0;
  assign cparam_matmul_33_out_col_step = 20;
  assign cparam_matmul_33_out_row_step = 20;
  assign cparam_matmul_33_out_bat_step = 20;
  assign cparam_matmul_33_out_och_step = 4;
  assign cparam_matmul_33_out_write_size = 1;
  assign cparam_matmul_33_out_write_size_res = 1;
  assign cparam_matmul_33_out_write_block = 0;
  assign cparam_matmul_33_keep_filter = 0;
  assign cparam_matmul_33_keep_input = 1;
  assign cparam_matmul_33_data_stationary = 0;
  assign cparam_matmul_33_stream_num_ops = 1;
  assign cparam_matmul_33_stream_num_ops_res = 1;
  assign cparam_matmul_33_stream_num_ops_par = 1;
  assign cparam_matmul_33_stream_num_ops_res_par = 1;
  assign cparam_matmul_33_stream_reduce_size = 256;
  assign cparam_matmul_33_stream_aligned_reduce_size = 256;
  assign cparam_matmul_33_stream_omit_mask = 0;
  assign cparam_matmul_33_col_select_initval = 0;
  assign cparam_matmul_33_stride_col_par_col = 1;
  assign cparam_matmul_33_stride_row_par_row = 1;
  assign cparam_matmul_33_stride_col_mod_filter_num = 0;
  assign cparam_matmul_33_filter_num_col_minus_stride_col_mod = 1;
  assign cparam_matmul_33_inc_act_laddr_conds_0 = 0;
  assign cparam_matmul_33_inc_act_laddr_small = 256;
  assign cparam_matmul_33_inc_act_laddr_large = 256;
  assign cparam_matmul_33_inc_out_laddr_col = 5;
  assign cparam_matmul_33_stream_act_local_small_offset = 0;
  assign cparam_matmul_33_stream_act_local_large_offset = 0;
  assign cparam_matmul_33_stream_act_local_small_flags_0 = 0;
  assign cparam_matmul_33_stream_act_local_large_flags_0 = 0;
  assign cparam_matmul_33_inc_sync_out = 1;
  assign cparam_matmul_33_inc_sync_out_res = 0;
  reg _acc_0_stream_ivalid;
  wire _acc_0_stream_oready;
  wire _acc_0_stream_internal_oready;
  assign _acc_0_stream_internal_oready = 1;
  reg [32-1:0] _acc_0_fsm;
  localparam _acc_0_fsm_init = 0;
  wire _acc_0_run_flag;
  assign _acc_0_run_flag = 0;
  reg _acc_0_source_start;
  wire _acc_0_source_stop;
  reg _acc_0_source_busy;
  wire _acc_0_sink_start;
  wire _acc_0_sink_stop;
  wire _acc_0_sink_busy;
  wire _acc_0_busy;
  reg _acc_0_busy_reg;
  wire _acc_0_is_root;
  reg _acc_0_x_idle;
  reg [33-1:0] _acc_0_x_source_count;
  reg [5-1:0] _acc_0_x_source_mode;
  reg [16-1:0] _acc_0_x_source_generator_id;
  reg [32-1:0] _acc_0_x_source_offset;
  reg [33-1:0] _acc_0_x_source_size;
  reg [32-1:0] _acc_0_x_source_stride;
  reg [32-1:0] _acc_0_x_source_offset_buf;
  reg [33-1:0] _acc_0_x_source_size_buf;
  reg [32-1:0] _acc_0_x_source_stride_buf;
  reg [8-1:0] _acc_0_x_source_sel;
  reg [32-1:0] _acc_0_x_source_ram_raddr;
  reg _acc_0_x_source_ram_renable;
  wire [64-1:0] _acc_0_x_source_ram_rdata;
  reg _acc_0_x_source_fifo_deq;
  wire [64-1:0] _acc_0_x_source_fifo_rdata;
  reg [64-1:0] _acc_0_x_source_empty_data;
  reg _acc_0_rshift_idle;
  reg [33-1:0] _acc_0_rshift_source_count;
  reg [5-1:0] _acc_0_rshift_source_mode;
  reg [16-1:0] _acc_0_rshift_source_generator_id;
  reg [32-1:0] _acc_0_rshift_source_offset;
  reg [33-1:0] _acc_0_rshift_source_size;
  reg [32-1:0] _acc_0_rshift_source_stride;
  reg [32-1:0] _acc_0_rshift_source_offset_buf;
  reg [33-1:0] _acc_0_rshift_source_size_buf;
  reg [32-1:0] _acc_0_rshift_source_stride_buf;
  reg [8-1:0] _acc_0_rshift_source_sel;
  reg [32-1:0] _acc_0_rshift_source_ram_raddr;
  reg _acc_0_rshift_source_ram_renable;
  wire [32-1:0] _acc_0_rshift_source_ram_rdata;
  reg _acc_0_rshift_source_fifo_deq;
  wire [32-1:0] _acc_0_rshift_source_fifo_rdata;
  reg [32-1:0] _acc_0_rshift_source_empty_data;
  reg [32-1:0] _acc_0_size_next_parameter_data;
  reg [33-1:0] _acc_0_sum_sink_count;
  reg [5-1:0] _acc_0_sum_sink_mode;
  reg [16-1:0] _acc_0_sum_sink_generator_id;
  reg [32-1:0] _acc_0_sum_sink_offset;
  reg [33-1:0] _acc_0_sum_sink_size;
  reg [32-1:0] _acc_0_sum_sink_stride;
  reg [32-1:0] _acc_0_sum_sink_offset_buf;
  reg [33-1:0] _acc_0_sum_sink_size_buf;
  reg [32-1:0] _acc_0_sum_sink_stride_buf;
  reg [8-1:0] _acc_0_sum_sink_sel;
  reg [32-1:0] _acc_0_sum_sink_waddr;
  reg _acc_0_sum_sink_wenable;
  reg [64-1:0] _acc_0_sum_sink_wdata;
  reg _acc_0_sum_sink_fifo_enq;
  reg [64-1:0] _acc_0_sum_sink_fifo_wdata;
  reg [64-1:0] _acc_0_sum_sink_immediate;
  reg [33-1:0] _acc_0_valid_sink_count;
  reg [5-1:0] _acc_0_valid_sink_mode;
  reg [16-1:0] _acc_0_valid_sink_generator_id;
  reg [32-1:0] _acc_0_valid_sink_offset;
  reg [33-1:0] _acc_0_valid_sink_size;
  reg [32-1:0] _acc_0_valid_sink_stride;
  reg [32-1:0] _acc_0_valid_sink_offset_buf;
  reg [33-1:0] _acc_0_valid_sink_size_buf;
  reg [32-1:0] _acc_0_valid_sink_stride_buf;
  reg [8-1:0] _acc_0_valid_sink_sel;
  reg [32-1:0] _acc_0_valid_sink_waddr;
  reg _acc_0_valid_sink_wenable;
  reg [1-1:0] _acc_0_valid_sink_wdata;
  reg _acc_0_valid_sink_fifo_enq;
  reg [1-1:0] _acc_0_valid_sink_fifo_wdata;
  reg [1-1:0] _acc_0_valid_sink_immediate;
  reg _acc_1_stream_ivalid;
  wire _acc_1_stream_oready;
  wire _acc_1_stream_internal_oready;
  assign _acc_1_stream_internal_oready = 1;
  reg [32-1:0] _acc_1_fsm;
  localparam _acc_1_fsm_init = 0;
  wire _acc_1_run_flag;
  assign _acc_1_run_flag = 0;
  reg _acc_1_source_start;
  wire _acc_1_source_stop;
  reg _acc_1_source_busy;
  wire _acc_1_sink_start;
  wire _acc_1_sink_stop;
  wire _acc_1_sink_busy;
  wire _acc_1_busy;
  reg _acc_1_busy_reg;
  wire _acc_1_is_root;
  reg _acc_1_x_idle;
  reg [33-1:0] _acc_1_x_source_count;
  reg [5-1:0] _acc_1_x_source_mode;
  reg [16-1:0] _acc_1_x_source_generator_id;
  reg [32-1:0] _acc_1_x_source_offset;
  reg [33-1:0] _acc_1_x_source_size;
  reg [32-1:0] _acc_1_x_source_stride;
  reg [32-1:0] _acc_1_x_source_offset_buf;
  reg [33-1:0] _acc_1_x_source_size_buf;
  reg [32-1:0] _acc_1_x_source_stride_buf;
  reg [8-1:0] _acc_1_x_source_sel;
  reg [32-1:0] _acc_1_x_source_ram_raddr;
  reg _acc_1_x_source_ram_renable;
  wire [64-1:0] _acc_1_x_source_ram_rdata;
  reg _acc_1_x_source_fifo_deq;
  wire [64-1:0] _acc_1_x_source_fifo_rdata;
  reg [64-1:0] _acc_1_x_source_empty_data;
  reg _acc_1_rshift_idle;
  reg [33-1:0] _acc_1_rshift_source_count;
  reg [5-1:0] _acc_1_rshift_source_mode;
  reg [16-1:0] _acc_1_rshift_source_generator_id;
  reg [32-1:0] _acc_1_rshift_source_offset;
  reg [33-1:0] _acc_1_rshift_source_size;
  reg [32-1:0] _acc_1_rshift_source_stride;
  reg [32-1:0] _acc_1_rshift_source_offset_buf;
  reg [33-1:0] _acc_1_rshift_source_size_buf;
  reg [32-1:0] _acc_1_rshift_source_stride_buf;
  reg [8-1:0] _acc_1_rshift_source_sel;
  reg [32-1:0] _acc_1_rshift_source_ram_raddr;
  reg _acc_1_rshift_source_ram_renable;
  wire [32-1:0] _acc_1_rshift_source_ram_rdata;
  reg _acc_1_rshift_source_fifo_deq;
  wire [32-1:0] _acc_1_rshift_source_fifo_rdata;
  reg [32-1:0] _acc_1_rshift_source_empty_data;
  reg [32-1:0] _acc_1_size_next_parameter_data;
  reg [33-1:0] _acc_1_sum_sink_count;
  reg [5-1:0] _acc_1_sum_sink_mode;
  reg [16-1:0] _acc_1_sum_sink_generator_id;
  reg [32-1:0] _acc_1_sum_sink_offset;
  reg [33-1:0] _acc_1_sum_sink_size;
  reg [32-1:0] _acc_1_sum_sink_stride;
  reg [32-1:0] _acc_1_sum_sink_offset_buf;
  reg [33-1:0] _acc_1_sum_sink_size_buf;
  reg [32-1:0] _acc_1_sum_sink_stride_buf;
  reg [8-1:0] _acc_1_sum_sink_sel;
  reg [32-1:0] _acc_1_sum_sink_waddr;
  reg _acc_1_sum_sink_wenable;
  reg [64-1:0] _acc_1_sum_sink_wdata;
  reg _acc_1_sum_sink_fifo_enq;
  reg [64-1:0] _acc_1_sum_sink_fifo_wdata;
  reg [64-1:0] _acc_1_sum_sink_immediate;
  reg [33-1:0] _acc_1_valid_sink_count;
  reg [5-1:0] _acc_1_valid_sink_mode;
  reg [16-1:0] _acc_1_valid_sink_generator_id;
  reg [32-1:0] _acc_1_valid_sink_offset;
  reg [33-1:0] _acc_1_valid_sink_size;
  reg [32-1:0] _acc_1_valid_sink_stride;
  reg [32-1:0] _acc_1_valid_sink_offset_buf;
  reg [33-1:0] _acc_1_valid_sink_size_buf;
  reg [32-1:0] _acc_1_valid_sink_stride_buf;
  reg [8-1:0] _acc_1_valid_sink_sel;
  reg [32-1:0] _acc_1_valid_sink_waddr;
  reg _acc_1_valid_sink_wenable;
  reg [1-1:0] _acc_1_valid_sink_wdata;
  reg _acc_1_valid_sink_fifo_enq;
  reg [1-1:0] _acc_1_valid_sink_fifo_wdata;
  reg [1-1:0] _acc_1_valid_sink_immediate;
  reg _add_tree_2_stream_ivalid;
  wire _add_tree_2_stream_oready;
  wire _add_tree_2_stream_internal_oready;
  assign _add_tree_2_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_2_fsm;
  localparam _add_tree_2_fsm_init = 0;
  wire _add_tree_2_run_flag;
  assign _add_tree_2_run_flag = 0;
  reg _add_tree_2_source_start;
  wire _add_tree_2_source_stop;
  reg _add_tree_2_source_busy;
  wire _add_tree_2_sink_start;
  wire _add_tree_2_sink_stop;
  wire _add_tree_2_sink_busy;
  wire _add_tree_2_busy;
  reg _add_tree_2_busy_reg;
  wire _add_tree_2_is_root;
  reg _add_tree_2_var0_idle;
  reg [33-1:0] _add_tree_2_var0_source_count;
  reg [5-1:0] _add_tree_2_var0_source_mode;
  reg [16-1:0] _add_tree_2_var0_source_generator_id;
  reg [32-1:0] _add_tree_2_var0_source_offset;
  reg [33-1:0] _add_tree_2_var0_source_size;
  reg [32-1:0] _add_tree_2_var0_source_stride;
  reg [32-1:0] _add_tree_2_var0_source_offset_buf;
  reg [33-1:0] _add_tree_2_var0_source_size_buf;
  reg [32-1:0] _add_tree_2_var0_source_stride_buf;
  reg [8-1:0] _add_tree_2_var0_source_sel;
  reg [32-1:0] _add_tree_2_var0_source_ram_raddr;
  reg _add_tree_2_var0_source_ram_renable;
  wire [64-1:0] _add_tree_2_var0_source_ram_rdata;
  reg _add_tree_2_var0_source_fifo_deq;
  wire [64-1:0] _add_tree_2_var0_source_fifo_rdata;
  reg [64-1:0] _add_tree_2_var0_source_empty_data;
  reg [33-1:0] _add_tree_2_sum_sink_count;
  reg [5-1:0] _add_tree_2_sum_sink_mode;
  reg [16-1:0] _add_tree_2_sum_sink_generator_id;
  reg [32-1:0] _add_tree_2_sum_sink_offset;
  reg [33-1:0] _add_tree_2_sum_sink_size;
  reg [32-1:0] _add_tree_2_sum_sink_stride;
  reg [32-1:0] _add_tree_2_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_2_sum_sink_size_buf;
  reg [32-1:0] _add_tree_2_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_2_sum_sink_sel;
  reg [32-1:0] _add_tree_2_sum_sink_waddr;
  reg _add_tree_2_sum_sink_wenable;
  reg [64-1:0] _add_tree_2_sum_sink_wdata;
  reg _add_tree_2_sum_sink_fifo_enq;
  reg [64-1:0] _add_tree_2_sum_sink_fifo_wdata;
  reg [64-1:0] _add_tree_2_sum_sink_immediate;
  reg _add_tree_3_stream_ivalid;
  wire _add_tree_3_stream_oready;
  wire _add_tree_3_stream_internal_oready;
  assign _add_tree_3_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_3_fsm;
  localparam _add_tree_3_fsm_init = 0;
  wire _add_tree_3_run_flag;
  assign _add_tree_3_run_flag = 0;
  reg _add_tree_3_source_start;
  wire _add_tree_3_source_stop;
  reg _add_tree_3_source_busy;
  wire _add_tree_3_sink_start;
  wire _add_tree_3_sink_stop;
  wire _add_tree_3_sink_busy;
  wire _add_tree_3_busy;
  reg _add_tree_3_busy_reg;
  wire _add_tree_3_is_root;
  reg _add_tree_3_var0_idle;
  reg [33-1:0] _add_tree_3_var0_source_count;
  reg [5-1:0] _add_tree_3_var0_source_mode;
  reg [16-1:0] _add_tree_3_var0_source_generator_id;
  reg [32-1:0] _add_tree_3_var0_source_offset;
  reg [33-1:0] _add_tree_3_var0_source_size;
  reg [32-1:0] _add_tree_3_var0_source_stride;
  reg [32-1:0] _add_tree_3_var0_source_offset_buf;
  reg [33-1:0] _add_tree_3_var0_source_size_buf;
  reg [32-1:0] _add_tree_3_var0_source_stride_buf;
  reg [8-1:0] _add_tree_3_var0_source_sel;
  reg [32-1:0] _add_tree_3_var0_source_ram_raddr;
  reg _add_tree_3_var0_source_ram_renable;
  wire [64-1:0] _add_tree_3_var0_source_ram_rdata;
  reg _add_tree_3_var0_source_fifo_deq;
  wire [64-1:0] _add_tree_3_var0_source_fifo_rdata;
  reg [64-1:0] _add_tree_3_var0_source_empty_data;
  reg _add_tree_3_var1_idle;
  reg [33-1:0] _add_tree_3_var1_source_count;
  reg [5-1:0] _add_tree_3_var1_source_mode;
  reg [16-1:0] _add_tree_3_var1_source_generator_id;
  reg [32-1:0] _add_tree_3_var1_source_offset;
  reg [33-1:0] _add_tree_3_var1_source_size;
  reg [32-1:0] _add_tree_3_var1_source_stride;
  reg [32-1:0] _add_tree_3_var1_source_offset_buf;
  reg [33-1:0] _add_tree_3_var1_source_size_buf;
  reg [32-1:0] _add_tree_3_var1_source_stride_buf;
  reg [8-1:0] _add_tree_3_var1_source_sel;
  reg [32-1:0] _add_tree_3_var1_source_ram_raddr;
  reg _add_tree_3_var1_source_ram_renable;
  wire [64-1:0] _add_tree_3_var1_source_ram_rdata;
  reg _add_tree_3_var1_source_fifo_deq;
  wire [64-1:0] _add_tree_3_var1_source_fifo_rdata;
  reg [64-1:0] _add_tree_3_var1_source_empty_data;
  reg [33-1:0] _add_tree_3_sum_sink_count;
  reg [5-1:0] _add_tree_3_sum_sink_mode;
  reg [16-1:0] _add_tree_3_sum_sink_generator_id;
  reg [32-1:0] _add_tree_3_sum_sink_offset;
  reg [33-1:0] _add_tree_3_sum_sink_size;
  reg [32-1:0] _add_tree_3_sum_sink_stride;
  reg [32-1:0] _add_tree_3_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_3_sum_sink_size_buf;
  reg [32-1:0] _add_tree_3_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_3_sum_sink_sel;
  reg [32-1:0] _add_tree_3_sum_sink_waddr;
  reg _add_tree_3_sum_sink_wenable;
  reg [64-1:0] _add_tree_3_sum_sink_wdata;
  reg _add_tree_3_sum_sink_fifo_enq;
  reg [64-1:0] _add_tree_3_sum_sink_fifo_wdata;
  reg [64-1:0] _add_tree_3_sum_sink_immediate;
  reg _add_tree_4_stream_ivalid;
  wire _add_tree_4_stream_oready;
  wire _add_tree_4_stream_internal_oready;
  assign _add_tree_4_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_4_fsm;
  localparam _add_tree_4_fsm_init = 0;
  wire _add_tree_4_run_flag;
  assign _add_tree_4_run_flag = 0;
  reg _add_tree_4_source_start;
  wire _add_tree_4_source_stop;
  reg _add_tree_4_source_busy;
  wire _add_tree_4_sink_start;
  wire _add_tree_4_sink_stop;
  wire _add_tree_4_sink_busy;
  wire _add_tree_4_busy;
  reg _add_tree_4_busy_reg;
  wire _add_tree_4_is_root;
  reg _add_tree_4_var0_idle;
  reg [33-1:0] _add_tree_4_var0_source_count;
  reg [5-1:0] _add_tree_4_var0_source_mode;
  reg [16-1:0] _add_tree_4_var0_source_generator_id;
  reg [32-1:0] _add_tree_4_var0_source_offset;
  reg [33-1:0] _add_tree_4_var0_source_size;
  reg [32-1:0] _add_tree_4_var0_source_stride;
  reg [32-1:0] _add_tree_4_var0_source_offset_buf;
  reg [33-1:0] _add_tree_4_var0_source_size_buf;
  reg [32-1:0] _add_tree_4_var0_source_stride_buf;
  reg [8-1:0] _add_tree_4_var0_source_sel;
  reg [32-1:0] _add_tree_4_var0_source_ram_raddr;
  reg _add_tree_4_var0_source_ram_renable;
  wire [64-1:0] _add_tree_4_var0_source_ram_rdata;
  reg _add_tree_4_var0_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var0_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var0_source_empty_data;
  reg _add_tree_4_var1_idle;
  reg [33-1:0] _add_tree_4_var1_source_count;
  reg [5-1:0] _add_tree_4_var1_source_mode;
  reg [16-1:0] _add_tree_4_var1_source_generator_id;
  reg [32-1:0] _add_tree_4_var1_source_offset;
  reg [33-1:0] _add_tree_4_var1_source_size;
  reg [32-1:0] _add_tree_4_var1_source_stride;
  reg [32-1:0] _add_tree_4_var1_source_offset_buf;
  reg [33-1:0] _add_tree_4_var1_source_size_buf;
  reg [32-1:0] _add_tree_4_var1_source_stride_buf;
  reg [8-1:0] _add_tree_4_var1_source_sel;
  reg [32-1:0] _add_tree_4_var1_source_ram_raddr;
  reg _add_tree_4_var1_source_ram_renable;
  wire [64-1:0] _add_tree_4_var1_source_ram_rdata;
  reg _add_tree_4_var1_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var1_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var1_source_empty_data;
  reg [33-1:0] _add_tree_4_sum_sink_count;
  reg [5-1:0] _add_tree_4_sum_sink_mode;
  reg [16-1:0] _add_tree_4_sum_sink_generator_id;
  reg [32-1:0] _add_tree_4_sum_sink_offset;
  reg [33-1:0] _add_tree_4_sum_sink_size;
  reg [32-1:0] _add_tree_4_sum_sink_stride;
  reg [32-1:0] _add_tree_4_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_4_sum_sink_size_buf;
  reg [32-1:0] _add_tree_4_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_4_sum_sink_sel;
  reg [32-1:0] _add_tree_4_sum_sink_waddr;
  reg _add_tree_4_sum_sink_wenable;
  reg [64-1:0] _add_tree_4_sum_sink_wdata;
  reg _add_tree_4_sum_sink_fifo_enq;
  reg [64-1:0] _add_tree_4_sum_sink_fifo_wdata;
  reg [64-1:0] _add_tree_4_sum_sink_immediate;
  reg _add_tree_5_stream_ivalid;
  wire _add_tree_5_stream_oready;
  wire _add_tree_5_stream_internal_oready;
  assign _add_tree_5_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_5_fsm;
  localparam _add_tree_5_fsm_init = 0;
  wire _add_tree_5_run_flag;
  assign _add_tree_5_run_flag = 0;
  reg _add_tree_5_source_start;
  wire _add_tree_5_source_stop;
  reg _add_tree_5_source_busy;
  wire _add_tree_5_sink_start;
  wire _add_tree_5_sink_stop;
  wire _add_tree_5_sink_busy;
  wire _add_tree_5_busy;
  reg _add_tree_5_busy_reg;
  wire _add_tree_5_is_root;
  reg _add_tree_5_var0_idle;
  reg [33-1:0] _add_tree_5_var0_source_count;
  reg [5-1:0] _add_tree_5_var0_source_mode;
  reg [16-1:0] _add_tree_5_var0_source_generator_id;
  reg [32-1:0] _add_tree_5_var0_source_offset;
  reg [33-1:0] _add_tree_5_var0_source_size;
  reg [32-1:0] _add_tree_5_var0_source_stride;
  reg [32-1:0] _add_tree_5_var0_source_offset_buf;
  reg [33-1:0] _add_tree_5_var0_source_size_buf;
  reg [32-1:0] _add_tree_5_var0_source_stride_buf;
  reg [8-1:0] _add_tree_5_var0_source_sel;
  reg [32-1:0] _add_tree_5_var0_source_ram_raddr;
  reg _add_tree_5_var0_source_ram_renable;
  wire [64-1:0] _add_tree_5_var0_source_ram_rdata;
  reg _add_tree_5_var0_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var0_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var0_source_empty_data;
  reg _add_tree_5_var1_idle;
  reg [33-1:0] _add_tree_5_var1_source_count;
  reg [5-1:0] _add_tree_5_var1_source_mode;
  reg [16-1:0] _add_tree_5_var1_source_generator_id;
  reg [32-1:0] _add_tree_5_var1_source_offset;
  reg [33-1:0] _add_tree_5_var1_source_size;
  reg [32-1:0] _add_tree_5_var1_source_stride;
  reg [32-1:0] _add_tree_5_var1_source_offset_buf;
  reg [33-1:0] _add_tree_5_var1_source_size_buf;
  reg [32-1:0] _add_tree_5_var1_source_stride_buf;
  reg [8-1:0] _add_tree_5_var1_source_sel;
  reg [32-1:0] _add_tree_5_var1_source_ram_raddr;
  reg _add_tree_5_var1_source_ram_renable;
  wire [64-1:0] _add_tree_5_var1_source_ram_rdata;
  reg _add_tree_5_var1_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var1_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var1_source_empty_data;
  reg _add_tree_5_var2_idle;
  reg [33-1:0] _add_tree_5_var2_source_count;
  reg [5-1:0] _add_tree_5_var2_source_mode;
  reg [16-1:0] _add_tree_5_var2_source_generator_id;
  reg [32-1:0] _add_tree_5_var2_source_offset;
  reg [33-1:0] _add_tree_5_var2_source_size;
  reg [32-1:0] _add_tree_5_var2_source_stride;
  reg [32-1:0] _add_tree_5_var2_source_offset_buf;
  reg [33-1:0] _add_tree_5_var2_source_size_buf;
  reg [32-1:0] _add_tree_5_var2_source_stride_buf;
  reg [8-1:0] _add_tree_5_var2_source_sel;
  reg [32-1:0] _add_tree_5_var2_source_ram_raddr;
  reg _add_tree_5_var2_source_ram_renable;
  wire [64-1:0] _add_tree_5_var2_source_ram_rdata;
  reg _add_tree_5_var2_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var2_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var2_source_empty_data;
  reg _add_tree_5_var3_idle;
  reg [33-1:0] _add_tree_5_var3_source_count;
  reg [5-1:0] _add_tree_5_var3_source_mode;
  reg [16-1:0] _add_tree_5_var3_source_generator_id;
  reg [32-1:0] _add_tree_5_var3_source_offset;
  reg [33-1:0] _add_tree_5_var3_source_size;
  reg [32-1:0] _add_tree_5_var3_source_stride;
  reg [32-1:0] _add_tree_5_var3_source_offset_buf;
  reg [33-1:0] _add_tree_5_var3_source_size_buf;
  reg [32-1:0] _add_tree_5_var3_source_stride_buf;
  reg [8-1:0] _add_tree_5_var3_source_sel;
  reg [32-1:0] _add_tree_5_var3_source_ram_raddr;
  reg _add_tree_5_var3_source_ram_renable;
  wire [64-1:0] _add_tree_5_var3_source_ram_rdata;
  reg _add_tree_5_var3_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var3_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var3_source_empty_data;
  reg _add_tree_5_var4_idle;
  reg [33-1:0] _add_tree_5_var4_source_count;
  reg [5-1:0] _add_tree_5_var4_source_mode;
  reg [16-1:0] _add_tree_5_var4_source_generator_id;
  reg [32-1:0] _add_tree_5_var4_source_offset;
  reg [33-1:0] _add_tree_5_var4_source_size;
  reg [32-1:0] _add_tree_5_var4_source_stride;
  reg [32-1:0] _add_tree_5_var4_source_offset_buf;
  reg [33-1:0] _add_tree_5_var4_source_size_buf;
  reg [32-1:0] _add_tree_5_var4_source_stride_buf;
  reg [8-1:0] _add_tree_5_var4_source_sel;
  reg [32-1:0] _add_tree_5_var4_source_ram_raddr;
  reg _add_tree_5_var4_source_ram_renable;
  wire [64-1:0] _add_tree_5_var4_source_ram_rdata;
  reg _add_tree_5_var4_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var4_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var4_source_empty_data;
  reg _add_tree_5_var5_idle;
  reg [33-1:0] _add_tree_5_var5_source_count;
  reg [5-1:0] _add_tree_5_var5_source_mode;
  reg [16-1:0] _add_tree_5_var5_source_generator_id;
  reg [32-1:0] _add_tree_5_var5_source_offset;
  reg [33-1:0] _add_tree_5_var5_source_size;
  reg [32-1:0] _add_tree_5_var5_source_stride;
  reg [32-1:0] _add_tree_5_var5_source_offset_buf;
  reg [33-1:0] _add_tree_5_var5_source_size_buf;
  reg [32-1:0] _add_tree_5_var5_source_stride_buf;
  reg [8-1:0] _add_tree_5_var5_source_sel;
  reg [32-1:0] _add_tree_5_var5_source_ram_raddr;
  reg _add_tree_5_var5_source_ram_renable;
  wire [64-1:0] _add_tree_5_var5_source_ram_rdata;
  reg _add_tree_5_var5_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var5_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var5_source_empty_data;
  reg _add_tree_5_var6_idle;
  reg [33-1:0] _add_tree_5_var6_source_count;
  reg [5-1:0] _add_tree_5_var6_source_mode;
  reg [16-1:0] _add_tree_5_var6_source_generator_id;
  reg [32-1:0] _add_tree_5_var6_source_offset;
  reg [33-1:0] _add_tree_5_var6_source_size;
  reg [32-1:0] _add_tree_5_var6_source_stride;
  reg [32-1:0] _add_tree_5_var6_source_offset_buf;
  reg [33-1:0] _add_tree_5_var6_source_size_buf;
  reg [32-1:0] _add_tree_5_var6_source_stride_buf;
  reg [8-1:0] _add_tree_5_var6_source_sel;
  reg [32-1:0] _add_tree_5_var6_source_ram_raddr;
  reg _add_tree_5_var6_source_ram_renable;
  wire [64-1:0] _add_tree_5_var6_source_ram_rdata;
  reg _add_tree_5_var6_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var6_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var6_source_empty_data;
  reg _add_tree_5_var7_idle;
  reg [33-1:0] _add_tree_5_var7_source_count;
  reg [5-1:0] _add_tree_5_var7_source_mode;
  reg [16-1:0] _add_tree_5_var7_source_generator_id;
  reg [32-1:0] _add_tree_5_var7_source_offset;
  reg [33-1:0] _add_tree_5_var7_source_size;
  reg [32-1:0] _add_tree_5_var7_source_stride;
  reg [32-1:0] _add_tree_5_var7_source_offset_buf;
  reg [33-1:0] _add_tree_5_var7_source_size_buf;
  reg [32-1:0] _add_tree_5_var7_source_stride_buf;
  reg [8-1:0] _add_tree_5_var7_source_sel;
  reg [32-1:0] _add_tree_5_var7_source_ram_raddr;
  reg _add_tree_5_var7_source_ram_renable;
  wire [64-1:0] _add_tree_5_var7_source_ram_rdata;
  reg _add_tree_5_var7_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var7_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var7_source_empty_data;
  reg _add_tree_5_var8_idle;
  reg [33-1:0] _add_tree_5_var8_source_count;
  reg [5-1:0] _add_tree_5_var8_source_mode;
  reg [16-1:0] _add_tree_5_var8_source_generator_id;
  reg [32-1:0] _add_tree_5_var8_source_offset;
  reg [33-1:0] _add_tree_5_var8_source_size;
  reg [32-1:0] _add_tree_5_var8_source_stride;
  reg [32-1:0] _add_tree_5_var8_source_offset_buf;
  reg [33-1:0] _add_tree_5_var8_source_size_buf;
  reg [32-1:0] _add_tree_5_var8_source_stride_buf;
  reg [8-1:0] _add_tree_5_var8_source_sel;
  reg [32-1:0] _add_tree_5_var8_source_ram_raddr;
  reg _add_tree_5_var8_source_ram_renable;
  wire [64-1:0] _add_tree_5_var8_source_ram_rdata;
  reg _add_tree_5_var8_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var8_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var8_source_empty_data;
  reg [33-1:0] _add_tree_5_sum_sink_count;
  reg [5-1:0] _add_tree_5_sum_sink_mode;
  reg [16-1:0] _add_tree_5_sum_sink_generator_id;
  reg [32-1:0] _add_tree_5_sum_sink_offset;
  reg [33-1:0] _add_tree_5_sum_sink_size;
  reg [32-1:0] _add_tree_5_sum_sink_stride;
  reg [32-1:0] _add_tree_5_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_5_sum_sink_size_buf;
  reg [32-1:0] _add_tree_5_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_5_sum_sink_sel;
  reg [32-1:0] _add_tree_5_sum_sink_waddr;
  reg _add_tree_5_sum_sink_wenable;
  reg [64-1:0] _add_tree_5_sum_sink_wdata;
  reg _add_tree_5_sum_sink_fifo_enq;
  reg [64-1:0] _add_tree_5_sum_sink_fifo_wdata;
  reg [64-1:0] _add_tree_5_sum_sink_immediate;
  reg _mul_rshift_round_clip_6_stream_ivalid;
  wire _mul_rshift_round_clip_6_stream_oready;
  wire _mul_rshift_round_clip_6_stream_internal_oready;
  assign _mul_rshift_round_clip_6_stream_internal_oready = 1;
  reg [32-1:0] _mul_rshift_round_clip_6_fsm;
  localparam _mul_rshift_round_clip_6_fsm_init = 0;
  wire _mul_rshift_round_clip_6_run_flag;
  assign _mul_rshift_round_clip_6_run_flag = 0;
  reg _mul_rshift_round_clip_6_source_start;
  wire _mul_rshift_round_clip_6_source_stop;
  reg _mul_rshift_round_clip_6_source_busy;
  wire _mul_rshift_round_clip_6_sink_start;
  wire _mul_rshift_round_clip_6_sink_stop;
  wire _mul_rshift_round_clip_6_sink_busy;
  wire _mul_rshift_round_clip_6_busy;
  reg _mul_rshift_round_clip_6_busy_reg;
  wire _mul_rshift_round_clip_6_is_root;
  reg _mul_rshift_round_clip_6_x_idle;
  reg [33-1:0] _mul_rshift_round_clip_6_x_source_count;
  reg [5-1:0] _mul_rshift_round_clip_6_x_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_6_x_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_6_x_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_6_x_source_size;
  reg [32-1:0] _mul_rshift_round_clip_6_x_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_6_x_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_6_x_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_6_x_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_6_x_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_6_x_source_ram_raddr;
  reg _mul_rshift_round_clip_6_x_source_ram_renable;
  wire [64-1:0] _mul_rshift_round_clip_6_x_source_ram_rdata;
  reg _mul_rshift_round_clip_6_x_source_fifo_deq;
  wire [64-1:0] _mul_rshift_round_clip_6_x_source_fifo_rdata;
  reg [64-1:0] _mul_rshift_round_clip_6_x_source_empty_data;
  reg _mul_rshift_round_clip_6_y_idle;
  reg [33-1:0] _mul_rshift_round_clip_6_y_source_count;
  reg [5-1:0] _mul_rshift_round_clip_6_y_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_6_y_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_6_y_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_6_y_source_size;
  reg [32-1:0] _mul_rshift_round_clip_6_y_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_6_y_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_6_y_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_6_y_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_6_y_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_6_y_source_ram_raddr;
  reg _mul_rshift_round_clip_6_y_source_ram_renable;
  wire [16-1:0] _mul_rshift_round_clip_6_y_source_ram_rdata;
  reg _mul_rshift_round_clip_6_y_source_fifo_deq;
  wire [16-1:0] _mul_rshift_round_clip_6_y_source_fifo_rdata;
  reg [16-1:0] _mul_rshift_round_clip_6_y_source_empty_data;
  reg _mul_rshift_round_clip_6_rshift_idle;
  reg [33-1:0] _mul_rshift_round_clip_6_rshift_source_count;
  reg [5-1:0] _mul_rshift_round_clip_6_rshift_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_6_rshift_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_6_rshift_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_6_rshift_source_size;
  reg [32-1:0] _mul_rshift_round_clip_6_rshift_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_6_rshift_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_6_rshift_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_6_rshift_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_6_rshift_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_6_rshift_source_ram_raddr;
  reg _mul_rshift_round_clip_6_rshift_source_ram_renable;
  wire [32-1:0] _mul_rshift_round_clip_6_rshift_source_ram_rdata;
  reg _mul_rshift_round_clip_6_rshift_source_fifo_deq;
  wire [32-1:0] _mul_rshift_round_clip_6_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_rshift_round_clip_6_rshift_source_empty_data;
  reg [33-1:0] _mul_rshift_round_clip_6_z_sink_count;
  reg [5-1:0] _mul_rshift_round_clip_6_z_sink_mode;
  reg [16-1:0] _mul_rshift_round_clip_6_z_sink_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_6_z_sink_offset;
  reg [33-1:0] _mul_rshift_round_clip_6_z_sink_size;
  reg [32-1:0] _mul_rshift_round_clip_6_z_sink_stride;
  reg [32-1:0] _mul_rshift_round_clip_6_z_sink_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_6_z_sink_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_6_z_sink_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_6_z_sink_sel;
  reg [32-1:0] _mul_rshift_round_clip_6_z_sink_waddr;
  reg _mul_rshift_round_clip_6_z_sink_wenable;
  reg [16-1:0] _mul_rshift_round_clip_6_z_sink_wdata;
  reg _mul_rshift_round_clip_6_z_sink_fifo_enq;
  reg [16-1:0] _mul_rshift_round_clip_6_z_sink_fifo_wdata;
  reg [16-1:0] _mul_rshift_round_clip_6_z_sink_immediate;
  reg _mul_rshift_round_clip_7_stream_ivalid;
  wire _mul_rshift_round_clip_7_stream_oready;
  wire _mul_rshift_round_clip_7_stream_internal_oready;
  assign _mul_rshift_round_clip_7_stream_internal_oready = 1;
  reg [32-1:0] _mul_rshift_round_clip_7_fsm;
  localparam _mul_rshift_round_clip_7_fsm_init = 0;
  wire _mul_rshift_round_clip_7_run_flag;
  assign _mul_rshift_round_clip_7_run_flag = 0;
  reg _mul_rshift_round_clip_7_source_start;
  wire _mul_rshift_round_clip_7_source_stop;
  reg _mul_rshift_round_clip_7_source_busy;
  wire _mul_rshift_round_clip_7_sink_start;
  wire _mul_rshift_round_clip_7_sink_stop;
  wire _mul_rshift_round_clip_7_sink_busy;
  wire _mul_rshift_round_clip_7_busy;
  reg _mul_rshift_round_clip_7_busy_reg;
  wire _mul_rshift_round_clip_7_is_root;
  reg _mul_rshift_round_clip_7_x_idle;
  reg [33-1:0] _mul_rshift_round_clip_7_x_source_count;
  reg [5-1:0] _mul_rshift_round_clip_7_x_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_7_x_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_7_x_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_7_x_source_size;
  reg [32-1:0] _mul_rshift_round_clip_7_x_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_7_x_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_7_x_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_7_x_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_7_x_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_7_x_source_ram_raddr;
  reg _mul_rshift_round_clip_7_x_source_ram_renable;
  wire [64-1:0] _mul_rshift_round_clip_7_x_source_ram_rdata;
  reg _mul_rshift_round_clip_7_x_source_fifo_deq;
  wire [64-1:0] _mul_rshift_round_clip_7_x_source_fifo_rdata;
  reg [64-1:0] _mul_rshift_round_clip_7_x_source_empty_data;
  reg _mul_rshift_round_clip_7_y_idle;
  reg [33-1:0] _mul_rshift_round_clip_7_y_source_count;
  reg [5-1:0] _mul_rshift_round_clip_7_y_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_7_y_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_7_y_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_7_y_source_size;
  reg [32-1:0] _mul_rshift_round_clip_7_y_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_7_y_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_7_y_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_7_y_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_7_y_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_7_y_source_ram_raddr;
  reg _mul_rshift_round_clip_7_y_source_ram_renable;
  wire [16-1:0] _mul_rshift_round_clip_7_y_source_ram_rdata;
  reg _mul_rshift_round_clip_7_y_source_fifo_deq;
  wire [16-1:0] _mul_rshift_round_clip_7_y_source_fifo_rdata;
  reg [16-1:0] _mul_rshift_round_clip_7_y_source_empty_data;
  reg _mul_rshift_round_clip_7_rshift_idle;
  reg [33-1:0] _mul_rshift_round_clip_7_rshift_source_count;
  reg [5-1:0] _mul_rshift_round_clip_7_rshift_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_7_rshift_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_7_rshift_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_7_rshift_source_size;
  reg [32-1:0] _mul_rshift_round_clip_7_rshift_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_7_rshift_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_7_rshift_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_7_rshift_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_7_rshift_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_7_rshift_source_ram_raddr;
  reg _mul_rshift_round_clip_7_rshift_source_ram_renable;
  wire [32-1:0] _mul_rshift_round_clip_7_rshift_source_ram_rdata;
  reg _mul_rshift_round_clip_7_rshift_source_fifo_deq;
  wire [32-1:0] _mul_rshift_round_clip_7_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_rshift_round_clip_7_rshift_source_empty_data;
  reg [33-1:0] _mul_rshift_round_clip_7_z_sink_count;
  reg [5-1:0] _mul_rshift_round_clip_7_z_sink_mode;
  reg [16-1:0] _mul_rshift_round_clip_7_z_sink_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_7_z_sink_offset;
  reg [33-1:0] _mul_rshift_round_clip_7_z_sink_size;
  reg [32-1:0] _mul_rshift_round_clip_7_z_sink_stride;
  reg [32-1:0] _mul_rshift_round_clip_7_z_sink_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_7_z_sink_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_7_z_sink_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_7_z_sink_sel;
  reg [32-1:0] _mul_rshift_round_clip_7_z_sink_waddr;
  reg _mul_rshift_round_clip_7_z_sink_wenable;
  reg [16-1:0] _mul_rshift_round_clip_7_z_sink_wdata;
  reg _mul_rshift_round_clip_7_z_sink_fifo_enq;
  reg [16-1:0] _mul_rshift_round_clip_7_z_sink_fifo_wdata;
  reg [16-1:0] _mul_rshift_round_clip_7_z_sink_immediate;
  reg _mul_8_stream_ivalid;
  wire _mul_8_stream_oready;
  wire _mul_8_stream_internal_oready;
  assign _mul_8_stream_internal_oready = 1;
  reg [32-1:0] _mul_8_fsm;
  localparam _mul_8_fsm_init = 0;
  wire _mul_8_run_flag;
  assign _mul_8_run_flag = 0;
  reg _mul_8_source_start;
  wire _mul_8_source_stop;
  reg _mul_8_source_busy;
  wire _mul_8_sink_start;
  wire _mul_8_sink_stop;
  wire _mul_8_sink_busy;
  wire _mul_8_busy;
  reg _mul_8_busy_reg;
  wire _mul_8_is_root;
  reg _mul_8_x_idle;
  reg [33-1:0] _mul_8_x_source_count;
  reg [5-1:0] _mul_8_x_source_mode;
  reg [16-1:0] _mul_8_x_source_generator_id;
  reg [32-1:0] _mul_8_x_source_offset;
  reg [33-1:0] _mul_8_x_source_size;
  reg [32-1:0] _mul_8_x_source_stride;
  reg [32-1:0] _mul_8_x_source_offset_buf;
  reg [33-1:0] _mul_8_x_source_size_buf;
  reg [32-1:0] _mul_8_x_source_stride_buf;
  reg [8-1:0] _mul_8_x_source_sel;
  reg [32-1:0] _mul_8_x_source_ram_raddr;
  reg _mul_8_x_source_ram_renable;
  wire [16-1:0] _mul_8_x_source_ram_rdata;
  reg _mul_8_x_source_fifo_deq;
  wire [16-1:0] _mul_8_x_source_fifo_rdata;
  reg [16-1:0] _mul_8_x_source_empty_data;
  reg _mul_8_y_idle;
  reg [33-1:0] _mul_8_y_source_count;
  reg [5-1:0] _mul_8_y_source_mode;
  reg [16-1:0] _mul_8_y_source_generator_id;
  reg [32-1:0] _mul_8_y_source_offset;
  reg [33-1:0] _mul_8_y_source_size;
  reg [32-1:0] _mul_8_y_source_stride;
  reg [32-1:0] _mul_8_y_source_offset_buf;
  reg [33-1:0] _mul_8_y_source_size_buf;
  reg [32-1:0] _mul_8_y_source_stride_buf;
  reg [8-1:0] _mul_8_y_source_sel;
  reg [32-1:0] _mul_8_y_source_ram_raddr;
  reg _mul_8_y_source_ram_renable;
  wire [16-1:0] _mul_8_y_source_ram_rdata;
  reg _mul_8_y_source_fifo_deq;
  wire [16-1:0] _mul_8_y_source_fifo_rdata;
  reg [16-1:0] _mul_8_y_source_empty_data;
  reg _mul_8_rshift_idle;
  reg [33-1:0] _mul_8_rshift_source_count;
  reg [5-1:0] _mul_8_rshift_source_mode;
  reg [16-1:0] _mul_8_rshift_source_generator_id;
  reg [32-1:0] _mul_8_rshift_source_offset;
  reg [33-1:0] _mul_8_rshift_source_size;
  reg [32-1:0] _mul_8_rshift_source_stride;
  reg [32-1:0] _mul_8_rshift_source_offset_buf;
  reg [33-1:0] _mul_8_rshift_source_size_buf;
  reg [32-1:0] _mul_8_rshift_source_stride_buf;
  reg [8-1:0] _mul_8_rshift_source_sel;
  reg [32-1:0] _mul_8_rshift_source_ram_raddr;
  reg _mul_8_rshift_source_ram_renable;
  wire [32-1:0] _mul_8_rshift_source_ram_rdata;
  reg _mul_8_rshift_source_fifo_deq;
  wire [32-1:0] _mul_8_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_8_rshift_source_empty_data;
  reg [33-1:0] _mul_8_z_sink_count;
  reg [5-1:0] _mul_8_z_sink_mode;
  reg [16-1:0] _mul_8_z_sink_generator_id;
  reg [32-1:0] _mul_8_z_sink_offset;
  reg [33-1:0] _mul_8_z_sink_size;
  reg [32-1:0] _mul_8_z_sink_stride;
  reg [32-1:0] _mul_8_z_sink_offset_buf;
  reg [33-1:0] _mul_8_z_sink_size_buf;
  reg [32-1:0] _mul_8_z_sink_stride_buf;
  reg [8-1:0] _mul_8_z_sink_sel;
  reg [32-1:0] _mul_8_z_sink_waddr;
  reg _mul_8_z_sink_wenable;
  reg [32-1:0] _mul_8_z_sink_wdata;
  reg _mul_8_z_sink_fifo_enq;
  reg [32-1:0] _mul_8_z_sink_fifo_wdata;
  reg [32-1:0] _mul_8_z_sink_immediate;
  reg _mul_9_stream_ivalid;
  wire _mul_9_stream_oready;
  wire _mul_9_stream_internal_oready;
  assign _mul_9_stream_internal_oready = 1;
  reg [32-1:0] _mul_9_fsm;
  localparam _mul_9_fsm_init = 0;
  wire _mul_9_run_flag;
  assign _mul_9_run_flag = 0;
  reg _mul_9_source_start;
  wire _mul_9_source_stop;
  reg _mul_9_source_busy;
  wire _mul_9_sink_start;
  wire _mul_9_sink_stop;
  wire _mul_9_sink_busy;
  wire _mul_9_busy;
  reg _mul_9_busy_reg;
  wire _mul_9_is_root;
  reg _mul_9_x_idle;
  reg [33-1:0] _mul_9_x_source_count;
  reg [5-1:0] _mul_9_x_source_mode;
  reg [16-1:0] _mul_9_x_source_generator_id;
  reg [32-1:0] _mul_9_x_source_offset;
  reg [33-1:0] _mul_9_x_source_size;
  reg [32-1:0] _mul_9_x_source_stride;
  reg [32-1:0] _mul_9_x_source_offset_buf;
  reg [33-1:0] _mul_9_x_source_size_buf;
  reg [32-1:0] _mul_9_x_source_stride_buf;
  reg [8-1:0] _mul_9_x_source_sel;
  reg [32-1:0] _mul_9_x_source_ram_raddr;
  reg _mul_9_x_source_ram_renable;
  wire [16-1:0] _mul_9_x_source_ram_rdata;
  reg _mul_9_x_source_fifo_deq;
  wire [16-1:0] _mul_9_x_source_fifo_rdata;
  reg [16-1:0] _mul_9_x_source_empty_data;
  reg _mul_9_y_idle;
  reg [33-1:0] _mul_9_y_source_count;
  reg [5-1:0] _mul_9_y_source_mode;
  reg [16-1:0] _mul_9_y_source_generator_id;
  reg [32-1:0] _mul_9_y_source_offset;
  reg [33-1:0] _mul_9_y_source_size;
  reg [32-1:0] _mul_9_y_source_stride;
  reg [32-1:0] _mul_9_y_source_offset_buf;
  reg [33-1:0] _mul_9_y_source_size_buf;
  reg [32-1:0] _mul_9_y_source_stride_buf;
  reg [8-1:0] _mul_9_y_source_sel;
  reg [32-1:0] _mul_9_y_source_ram_raddr;
  reg _mul_9_y_source_ram_renable;
  wire [16-1:0] _mul_9_y_source_ram_rdata;
  reg _mul_9_y_source_fifo_deq;
  wire [16-1:0] _mul_9_y_source_fifo_rdata;
  reg [16-1:0] _mul_9_y_source_empty_data;
  reg _mul_9_rshift_idle;
  reg [33-1:0] _mul_9_rshift_source_count;
  reg [5-1:0] _mul_9_rshift_source_mode;
  reg [16-1:0] _mul_9_rshift_source_generator_id;
  reg [32-1:0] _mul_9_rshift_source_offset;
  reg [33-1:0] _mul_9_rshift_source_size;
  reg [32-1:0] _mul_9_rshift_source_stride;
  reg [32-1:0] _mul_9_rshift_source_offset_buf;
  reg [33-1:0] _mul_9_rshift_source_size_buf;
  reg [32-1:0] _mul_9_rshift_source_stride_buf;
  reg [8-1:0] _mul_9_rshift_source_sel;
  reg [32-1:0] _mul_9_rshift_source_ram_raddr;
  reg _mul_9_rshift_source_ram_renable;
  wire [32-1:0] _mul_9_rshift_source_ram_rdata;
  reg _mul_9_rshift_source_fifo_deq;
  wire [32-1:0] _mul_9_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_9_rshift_source_empty_data;
  reg [33-1:0] _mul_9_z_sink_count;
  reg [5-1:0] _mul_9_z_sink_mode;
  reg [16-1:0] _mul_9_z_sink_generator_id;
  reg [32-1:0] _mul_9_z_sink_offset;
  reg [33-1:0] _mul_9_z_sink_size;
  reg [32-1:0] _mul_9_z_sink_stride;
  reg [32-1:0] _mul_9_z_sink_offset_buf;
  reg [33-1:0] _mul_9_z_sink_size_buf;
  reg [32-1:0] _mul_9_z_sink_stride_buf;
  reg [8-1:0] _mul_9_z_sink_sel;
  reg [32-1:0] _mul_9_z_sink_waddr;
  reg _mul_9_z_sink_wenable;
  reg [32-1:0] _mul_9_z_sink_wdata;
  reg _mul_9_z_sink_fifo_enq;
  reg [32-1:0] _mul_9_z_sink_fifo_wdata;
  reg [32-1:0] _mul_9_z_sink_immediate;
  reg _mul_10_stream_ivalid;
  wire _mul_10_stream_oready;
  wire _mul_10_stream_internal_oready;
  assign _mul_10_stream_internal_oready = 1;
  reg [32-1:0] _mul_10_fsm;
  localparam _mul_10_fsm_init = 0;
  wire _mul_10_run_flag;
  assign _mul_10_run_flag = 0;
  reg _mul_10_source_start;
  wire _mul_10_source_stop;
  reg _mul_10_source_busy;
  wire _mul_10_sink_start;
  wire _mul_10_sink_stop;
  wire _mul_10_sink_busy;
  wire _mul_10_busy;
  reg _mul_10_busy_reg;
  wire _mul_10_is_root;
  reg _mul_10_x_idle;
  reg [33-1:0] _mul_10_x_source_count;
  reg [5-1:0] _mul_10_x_source_mode;
  reg [16-1:0] _mul_10_x_source_generator_id;
  reg [32-1:0] _mul_10_x_source_offset;
  reg [33-1:0] _mul_10_x_source_size;
  reg [32-1:0] _mul_10_x_source_stride;
  reg [32-1:0] _mul_10_x_source_offset_buf;
  reg [33-1:0] _mul_10_x_source_size_buf;
  reg [32-1:0] _mul_10_x_source_stride_buf;
  reg [8-1:0] _mul_10_x_source_sel;
  reg [32-1:0] _mul_10_x_source_ram_raddr;
  reg _mul_10_x_source_ram_renable;
  wire [16-1:0] _mul_10_x_source_ram_rdata;
  reg _mul_10_x_source_fifo_deq;
  wire [16-1:0] _mul_10_x_source_fifo_rdata;
  reg [16-1:0] _mul_10_x_source_empty_data;
  reg _mul_10_y_idle;
  reg [33-1:0] _mul_10_y_source_count;
  reg [5-1:0] _mul_10_y_source_mode;
  reg [16-1:0] _mul_10_y_source_generator_id;
  reg [32-1:0] _mul_10_y_source_offset;
  reg [33-1:0] _mul_10_y_source_size;
  reg [32-1:0] _mul_10_y_source_stride;
  reg [32-1:0] _mul_10_y_source_offset_buf;
  reg [33-1:0] _mul_10_y_source_size_buf;
  reg [32-1:0] _mul_10_y_source_stride_buf;
  reg [8-1:0] _mul_10_y_source_sel;
  reg [32-1:0] _mul_10_y_source_ram_raddr;
  reg _mul_10_y_source_ram_renable;
  wire [16-1:0] _mul_10_y_source_ram_rdata;
  reg _mul_10_y_source_fifo_deq;
  wire [16-1:0] _mul_10_y_source_fifo_rdata;
  reg [16-1:0] _mul_10_y_source_empty_data;
  reg _mul_10_rshift_idle;
  reg [33-1:0] _mul_10_rshift_source_count;
  reg [5-1:0] _mul_10_rshift_source_mode;
  reg [16-1:0] _mul_10_rshift_source_generator_id;
  reg [32-1:0] _mul_10_rshift_source_offset;
  reg [33-1:0] _mul_10_rshift_source_size;
  reg [32-1:0] _mul_10_rshift_source_stride;
  reg [32-1:0] _mul_10_rshift_source_offset_buf;
  reg [33-1:0] _mul_10_rshift_source_size_buf;
  reg [32-1:0] _mul_10_rshift_source_stride_buf;
  reg [8-1:0] _mul_10_rshift_source_sel;
  reg [32-1:0] _mul_10_rshift_source_ram_raddr;
  reg _mul_10_rshift_source_ram_renable;
  wire [32-1:0] _mul_10_rshift_source_ram_rdata;
  reg _mul_10_rshift_source_fifo_deq;
  wire [32-1:0] _mul_10_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_10_rshift_source_empty_data;
  reg [33-1:0] _mul_10_z_sink_count;
  reg [5-1:0] _mul_10_z_sink_mode;
  reg [16-1:0] _mul_10_z_sink_generator_id;
  reg [32-1:0] _mul_10_z_sink_offset;
  reg [33-1:0] _mul_10_z_sink_size;
  reg [32-1:0] _mul_10_z_sink_stride;
  reg [32-1:0] _mul_10_z_sink_offset_buf;
  reg [33-1:0] _mul_10_z_sink_size_buf;
  reg [32-1:0] _mul_10_z_sink_stride_buf;
  reg [8-1:0] _mul_10_z_sink_sel;
  reg [32-1:0] _mul_10_z_sink_waddr;
  reg _mul_10_z_sink_wenable;
  reg [32-1:0] _mul_10_z_sink_wdata;
  reg _mul_10_z_sink_fifo_enq;
  reg [32-1:0] _mul_10_z_sink_fifo_wdata;
  reg [32-1:0] _mul_10_z_sink_immediate;
  reg _mul_11_stream_ivalid;
  wire _mul_11_stream_oready;
  wire _mul_11_stream_internal_oready;
  assign _mul_11_stream_internal_oready = 1;
  reg [32-1:0] _mul_11_fsm;
  localparam _mul_11_fsm_init = 0;
  wire _mul_11_run_flag;
  assign _mul_11_run_flag = 0;
  reg _mul_11_source_start;
  wire _mul_11_source_stop;
  reg _mul_11_source_busy;
  wire _mul_11_sink_start;
  wire _mul_11_sink_stop;
  wire _mul_11_sink_busy;
  wire _mul_11_busy;
  reg _mul_11_busy_reg;
  wire _mul_11_is_root;
  reg _mul_11_x_idle;
  reg [33-1:0] _mul_11_x_source_count;
  reg [5-1:0] _mul_11_x_source_mode;
  reg [16-1:0] _mul_11_x_source_generator_id;
  reg [32-1:0] _mul_11_x_source_offset;
  reg [33-1:0] _mul_11_x_source_size;
  reg [32-1:0] _mul_11_x_source_stride;
  reg [32-1:0] _mul_11_x_source_offset_buf;
  reg [33-1:0] _mul_11_x_source_size_buf;
  reg [32-1:0] _mul_11_x_source_stride_buf;
  reg [8-1:0] _mul_11_x_source_sel;
  reg [32-1:0] _mul_11_x_source_ram_raddr;
  reg _mul_11_x_source_ram_renable;
  wire [16-1:0] _mul_11_x_source_ram_rdata;
  reg _mul_11_x_source_fifo_deq;
  wire [16-1:0] _mul_11_x_source_fifo_rdata;
  reg [16-1:0] _mul_11_x_source_empty_data;
  reg _mul_11_y_idle;
  reg [33-1:0] _mul_11_y_source_count;
  reg [5-1:0] _mul_11_y_source_mode;
  reg [16-1:0] _mul_11_y_source_generator_id;
  reg [32-1:0] _mul_11_y_source_offset;
  reg [33-1:0] _mul_11_y_source_size;
  reg [32-1:0] _mul_11_y_source_stride;
  reg [32-1:0] _mul_11_y_source_offset_buf;
  reg [33-1:0] _mul_11_y_source_size_buf;
  reg [32-1:0] _mul_11_y_source_stride_buf;
  reg [8-1:0] _mul_11_y_source_sel;
  reg [32-1:0] _mul_11_y_source_ram_raddr;
  reg _mul_11_y_source_ram_renable;
  wire [16-1:0] _mul_11_y_source_ram_rdata;
  reg _mul_11_y_source_fifo_deq;
  wire [16-1:0] _mul_11_y_source_fifo_rdata;
  reg [16-1:0] _mul_11_y_source_empty_data;
  reg _mul_11_rshift_idle;
  reg [33-1:0] _mul_11_rshift_source_count;
  reg [5-1:0] _mul_11_rshift_source_mode;
  reg [16-1:0] _mul_11_rshift_source_generator_id;
  reg [32-1:0] _mul_11_rshift_source_offset;
  reg [33-1:0] _mul_11_rshift_source_size;
  reg [32-1:0] _mul_11_rshift_source_stride;
  reg [32-1:0] _mul_11_rshift_source_offset_buf;
  reg [33-1:0] _mul_11_rshift_source_size_buf;
  reg [32-1:0] _mul_11_rshift_source_stride_buf;
  reg [8-1:0] _mul_11_rshift_source_sel;
  reg [32-1:0] _mul_11_rshift_source_ram_raddr;
  reg _mul_11_rshift_source_ram_renable;
  wire [32-1:0] _mul_11_rshift_source_ram_rdata;
  reg _mul_11_rshift_source_fifo_deq;
  wire [32-1:0] _mul_11_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_11_rshift_source_empty_data;
  reg [33-1:0] _mul_11_z_sink_count;
  reg [5-1:0] _mul_11_z_sink_mode;
  reg [16-1:0] _mul_11_z_sink_generator_id;
  reg [32-1:0] _mul_11_z_sink_offset;
  reg [33-1:0] _mul_11_z_sink_size;
  reg [32-1:0] _mul_11_z_sink_stride;
  reg [32-1:0] _mul_11_z_sink_offset_buf;
  reg [33-1:0] _mul_11_z_sink_size_buf;
  reg [32-1:0] _mul_11_z_sink_stride_buf;
  reg [8-1:0] _mul_11_z_sink_sel;
  reg [32-1:0] _mul_11_z_sink_waddr;
  reg _mul_11_z_sink_wenable;
  reg [32-1:0] _mul_11_z_sink_wdata;
  reg _mul_11_z_sink_fifo_enq;
  reg [32-1:0] _mul_11_z_sink_fifo_wdata;
  reg [32-1:0] _mul_11_z_sink_immediate;
  reg _mul_12_stream_ivalid;
  wire _mul_12_stream_oready;
  wire _mul_12_stream_internal_oready;
  assign _mul_12_stream_internal_oready = 1;
  reg [32-1:0] _mul_12_fsm;
  localparam _mul_12_fsm_init = 0;
  wire _mul_12_run_flag;
  assign _mul_12_run_flag = 0;
  reg _mul_12_source_start;
  wire _mul_12_source_stop;
  reg _mul_12_source_busy;
  wire _mul_12_sink_start;
  wire _mul_12_sink_stop;
  wire _mul_12_sink_busy;
  wire _mul_12_busy;
  reg _mul_12_busy_reg;
  wire _mul_12_is_root;
  reg _mul_12_x_idle;
  reg [33-1:0] _mul_12_x_source_count;
  reg [5-1:0] _mul_12_x_source_mode;
  reg [16-1:0] _mul_12_x_source_generator_id;
  reg [32-1:0] _mul_12_x_source_offset;
  reg [33-1:0] _mul_12_x_source_size;
  reg [32-1:0] _mul_12_x_source_stride;
  reg [32-1:0] _mul_12_x_source_offset_buf;
  reg [33-1:0] _mul_12_x_source_size_buf;
  reg [32-1:0] _mul_12_x_source_stride_buf;
  reg [8-1:0] _mul_12_x_source_sel;
  reg [32-1:0] _mul_12_x_source_ram_raddr;
  reg _mul_12_x_source_ram_renable;
  wire [16-1:0] _mul_12_x_source_ram_rdata;
  reg _mul_12_x_source_fifo_deq;
  wire [16-1:0] _mul_12_x_source_fifo_rdata;
  reg [16-1:0] _mul_12_x_source_empty_data;
  reg _mul_12_y_idle;
  reg [33-1:0] _mul_12_y_source_count;
  reg [5-1:0] _mul_12_y_source_mode;
  reg [16-1:0] _mul_12_y_source_generator_id;
  reg [32-1:0] _mul_12_y_source_offset;
  reg [33-1:0] _mul_12_y_source_size;
  reg [32-1:0] _mul_12_y_source_stride;
  reg [32-1:0] _mul_12_y_source_offset_buf;
  reg [33-1:0] _mul_12_y_source_size_buf;
  reg [32-1:0] _mul_12_y_source_stride_buf;
  reg [8-1:0] _mul_12_y_source_sel;
  reg [32-1:0] _mul_12_y_source_ram_raddr;
  reg _mul_12_y_source_ram_renable;
  wire [16-1:0] _mul_12_y_source_ram_rdata;
  reg _mul_12_y_source_fifo_deq;
  wire [16-1:0] _mul_12_y_source_fifo_rdata;
  reg [16-1:0] _mul_12_y_source_empty_data;
  reg _mul_12_rshift_idle;
  reg [33-1:0] _mul_12_rshift_source_count;
  reg [5-1:0] _mul_12_rshift_source_mode;
  reg [16-1:0] _mul_12_rshift_source_generator_id;
  reg [32-1:0] _mul_12_rshift_source_offset;
  reg [33-1:0] _mul_12_rshift_source_size;
  reg [32-1:0] _mul_12_rshift_source_stride;
  reg [32-1:0] _mul_12_rshift_source_offset_buf;
  reg [33-1:0] _mul_12_rshift_source_size_buf;
  reg [32-1:0] _mul_12_rshift_source_stride_buf;
  reg [8-1:0] _mul_12_rshift_source_sel;
  reg [32-1:0] _mul_12_rshift_source_ram_raddr;
  reg _mul_12_rshift_source_ram_renable;
  wire [32-1:0] _mul_12_rshift_source_ram_rdata;
  reg _mul_12_rshift_source_fifo_deq;
  wire [32-1:0] _mul_12_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_12_rshift_source_empty_data;
  reg [33-1:0] _mul_12_z_sink_count;
  reg [5-1:0] _mul_12_z_sink_mode;
  reg [16-1:0] _mul_12_z_sink_generator_id;
  reg [32-1:0] _mul_12_z_sink_offset;
  reg [33-1:0] _mul_12_z_sink_size;
  reg [32-1:0] _mul_12_z_sink_stride;
  reg [32-1:0] _mul_12_z_sink_offset_buf;
  reg [33-1:0] _mul_12_z_sink_size_buf;
  reg [32-1:0] _mul_12_z_sink_stride_buf;
  reg [8-1:0] _mul_12_z_sink_sel;
  reg [32-1:0] _mul_12_z_sink_waddr;
  reg _mul_12_z_sink_wenable;
  reg [32-1:0] _mul_12_z_sink_wdata;
  reg _mul_12_z_sink_fifo_enq;
  reg [32-1:0] _mul_12_z_sink_fifo_wdata;
  reg [32-1:0] _mul_12_z_sink_immediate;
  reg _mul_13_stream_ivalid;
  wire _mul_13_stream_oready;
  wire _mul_13_stream_internal_oready;
  assign _mul_13_stream_internal_oready = 1;
  reg [32-1:0] _mul_13_fsm;
  localparam _mul_13_fsm_init = 0;
  wire _mul_13_run_flag;
  assign _mul_13_run_flag = 0;
  reg _mul_13_source_start;
  wire _mul_13_source_stop;
  reg _mul_13_source_busy;
  wire _mul_13_sink_start;
  wire _mul_13_sink_stop;
  wire _mul_13_sink_busy;
  wire _mul_13_busy;
  reg _mul_13_busy_reg;
  wire _mul_13_is_root;
  reg _mul_13_x_idle;
  reg [33-1:0] _mul_13_x_source_count;
  reg [5-1:0] _mul_13_x_source_mode;
  reg [16-1:0] _mul_13_x_source_generator_id;
  reg [32-1:0] _mul_13_x_source_offset;
  reg [33-1:0] _mul_13_x_source_size;
  reg [32-1:0] _mul_13_x_source_stride;
  reg [32-1:0] _mul_13_x_source_offset_buf;
  reg [33-1:0] _mul_13_x_source_size_buf;
  reg [32-1:0] _mul_13_x_source_stride_buf;
  reg [8-1:0] _mul_13_x_source_sel;
  reg [32-1:0] _mul_13_x_source_ram_raddr;
  reg _mul_13_x_source_ram_renable;
  wire [16-1:0] _mul_13_x_source_ram_rdata;
  reg _mul_13_x_source_fifo_deq;
  wire [16-1:0] _mul_13_x_source_fifo_rdata;
  reg [16-1:0] _mul_13_x_source_empty_data;
  reg _mul_13_y_idle;
  reg [33-1:0] _mul_13_y_source_count;
  reg [5-1:0] _mul_13_y_source_mode;
  reg [16-1:0] _mul_13_y_source_generator_id;
  reg [32-1:0] _mul_13_y_source_offset;
  reg [33-1:0] _mul_13_y_source_size;
  reg [32-1:0] _mul_13_y_source_stride;
  reg [32-1:0] _mul_13_y_source_offset_buf;
  reg [33-1:0] _mul_13_y_source_size_buf;
  reg [32-1:0] _mul_13_y_source_stride_buf;
  reg [8-1:0] _mul_13_y_source_sel;
  reg [32-1:0] _mul_13_y_source_ram_raddr;
  reg _mul_13_y_source_ram_renable;
  wire [16-1:0] _mul_13_y_source_ram_rdata;
  reg _mul_13_y_source_fifo_deq;
  wire [16-1:0] _mul_13_y_source_fifo_rdata;
  reg [16-1:0] _mul_13_y_source_empty_data;
  reg _mul_13_rshift_idle;
  reg [33-1:0] _mul_13_rshift_source_count;
  reg [5-1:0] _mul_13_rshift_source_mode;
  reg [16-1:0] _mul_13_rshift_source_generator_id;
  reg [32-1:0] _mul_13_rshift_source_offset;
  reg [33-1:0] _mul_13_rshift_source_size;
  reg [32-1:0] _mul_13_rshift_source_stride;
  reg [32-1:0] _mul_13_rshift_source_offset_buf;
  reg [33-1:0] _mul_13_rshift_source_size_buf;
  reg [32-1:0] _mul_13_rshift_source_stride_buf;
  reg [8-1:0] _mul_13_rshift_source_sel;
  reg [32-1:0] _mul_13_rshift_source_ram_raddr;
  reg _mul_13_rshift_source_ram_renable;
  wire [32-1:0] _mul_13_rshift_source_ram_rdata;
  reg _mul_13_rshift_source_fifo_deq;
  wire [32-1:0] _mul_13_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_13_rshift_source_empty_data;
  reg [33-1:0] _mul_13_z_sink_count;
  reg [5-1:0] _mul_13_z_sink_mode;
  reg [16-1:0] _mul_13_z_sink_generator_id;
  reg [32-1:0] _mul_13_z_sink_offset;
  reg [33-1:0] _mul_13_z_sink_size;
  reg [32-1:0] _mul_13_z_sink_stride;
  reg [32-1:0] _mul_13_z_sink_offset_buf;
  reg [33-1:0] _mul_13_z_sink_size_buf;
  reg [32-1:0] _mul_13_z_sink_stride_buf;
  reg [8-1:0] _mul_13_z_sink_sel;
  reg [32-1:0] _mul_13_z_sink_waddr;
  reg _mul_13_z_sink_wenable;
  reg [32-1:0] _mul_13_z_sink_wdata;
  reg _mul_13_z_sink_fifo_enq;
  reg [32-1:0] _mul_13_z_sink_fifo_wdata;
  reg [32-1:0] _mul_13_z_sink_immediate;
  reg _mul_14_stream_ivalid;
  wire _mul_14_stream_oready;
  wire _mul_14_stream_internal_oready;
  assign _mul_14_stream_internal_oready = 1;
  reg [32-1:0] _mul_14_fsm;
  localparam _mul_14_fsm_init = 0;
  wire _mul_14_run_flag;
  assign _mul_14_run_flag = 0;
  reg _mul_14_source_start;
  wire _mul_14_source_stop;
  reg _mul_14_source_busy;
  wire _mul_14_sink_start;
  wire _mul_14_sink_stop;
  wire _mul_14_sink_busy;
  wire _mul_14_busy;
  reg _mul_14_busy_reg;
  wire _mul_14_is_root;
  reg _mul_14_x_idle;
  reg [33-1:0] _mul_14_x_source_count;
  reg [5-1:0] _mul_14_x_source_mode;
  reg [16-1:0] _mul_14_x_source_generator_id;
  reg [32-1:0] _mul_14_x_source_offset;
  reg [33-1:0] _mul_14_x_source_size;
  reg [32-1:0] _mul_14_x_source_stride;
  reg [32-1:0] _mul_14_x_source_offset_buf;
  reg [33-1:0] _mul_14_x_source_size_buf;
  reg [32-1:0] _mul_14_x_source_stride_buf;
  reg [8-1:0] _mul_14_x_source_sel;
  reg [32-1:0] _mul_14_x_source_ram_raddr;
  reg _mul_14_x_source_ram_renable;
  wire [16-1:0] _mul_14_x_source_ram_rdata;
  reg _mul_14_x_source_fifo_deq;
  wire [16-1:0] _mul_14_x_source_fifo_rdata;
  reg [16-1:0] _mul_14_x_source_empty_data;
  reg _mul_14_y_idle;
  reg [33-1:0] _mul_14_y_source_count;
  reg [5-1:0] _mul_14_y_source_mode;
  reg [16-1:0] _mul_14_y_source_generator_id;
  reg [32-1:0] _mul_14_y_source_offset;
  reg [33-1:0] _mul_14_y_source_size;
  reg [32-1:0] _mul_14_y_source_stride;
  reg [32-1:0] _mul_14_y_source_offset_buf;
  reg [33-1:0] _mul_14_y_source_size_buf;
  reg [32-1:0] _mul_14_y_source_stride_buf;
  reg [8-1:0] _mul_14_y_source_sel;
  reg [32-1:0] _mul_14_y_source_ram_raddr;
  reg _mul_14_y_source_ram_renable;
  wire [16-1:0] _mul_14_y_source_ram_rdata;
  reg _mul_14_y_source_fifo_deq;
  wire [16-1:0] _mul_14_y_source_fifo_rdata;
  reg [16-1:0] _mul_14_y_source_empty_data;
  reg _mul_14_rshift_idle;
  reg [33-1:0] _mul_14_rshift_source_count;
  reg [5-1:0] _mul_14_rshift_source_mode;
  reg [16-1:0] _mul_14_rshift_source_generator_id;
  reg [32-1:0] _mul_14_rshift_source_offset;
  reg [33-1:0] _mul_14_rshift_source_size;
  reg [32-1:0] _mul_14_rshift_source_stride;
  reg [32-1:0] _mul_14_rshift_source_offset_buf;
  reg [33-1:0] _mul_14_rshift_source_size_buf;
  reg [32-1:0] _mul_14_rshift_source_stride_buf;
  reg [8-1:0] _mul_14_rshift_source_sel;
  reg [32-1:0] _mul_14_rshift_source_ram_raddr;
  reg _mul_14_rshift_source_ram_renable;
  wire [32-1:0] _mul_14_rshift_source_ram_rdata;
  reg _mul_14_rshift_source_fifo_deq;
  wire [32-1:0] _mul_14_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_14_rshift_source_empty_data;
  reg [33-1:0] _mul_14_z_sink_count;
  reg [5-1:0] _mul_14_z_sink_mode;
  reg [16-1:0] _mul_14_z_sink_generator_id;
  reg [32-1:0] _mul_14_z_sink_offset;
  reg [33-1:0] _mul_14_z_sink_size;
  reg [32-1:0] _mul_14_z_sink_stride;
  reg [32-1:0] _mul_14_z_sink_offset_buf;
  reg [33-1:0] _mul_14_z_sink_size_buf;
  reg [32-1:0] _mul_14_z_sink_stride_buf;
  reg [8-1:0] _mul_14_z_sink_sel;
  reg [32-1:0] _mul_14_z_sink_waddr;
  reg _mul_14_z_sink_wenable;
  reg [32-1:0] _mul_14_z_sink_wdata;
  reg _mul_14_z_sink_fifo_enq;
  reg [32-1:0] _mul_14_z_sink_fifo_wdata;
  reg [32-1:0] _mul_14_z_sink_immediate;
  reg _mul_15_stream_ivalid;
  wire _mul_15_stream_oready;
  wire _mul_15_stream_internal_oready;
  assign _mul_15_stream_internal_oready = 1;
  reg [32-1:0] _mul_15_fsm;
  localparam _mul_15_fsm_init = 0;
  wire _mul_15_run_flag;
  assign _mul_15_run_flag = 0;
  reg _mul_15_source_start;
  wire _mul_15_source_stop;
  reg _mul_15_source_busy;
  wire _mul_15_sink_start;
  wire _mul_15_sink_stop;
  wire _mul_15_sink_busy;
  wire _mul_15_busy;
  reg _mul_15_busy_reg;
  wire _mul_15_is_root;
  reg _mul_15_x_idle;
  reg [33-1:0] _mul_15_x_source_count;
  reg [5-1:0] _mul_15_x_source_mode;
  reg [16-1:0] _mul_15_x_source_generator_id;
  reg [32-1:0] _mul_15_x_source_offset;
  reg [33-1:0] _mul_15_x_source_size;
  reg [32-1:0] _mul_15_x_source_stride;
  reg [32-1:0] _mul_15_x_source_offset_buf;
  reg [33-1:0] _mul_15_x_source_size_buf;
  reg [32-1:0] _mul_15_x_source_stride_buf;
  reg [8-1:0] _mul_15_x_source_sel;
  reg [32-1:0] _mul_15_x_source_ram_raddr;
  reg _mul_15_x_source_ram_renable;
  wire [16-1:0] _mul_15_x_source_ram_rdata;
  reg _mul_15_x_source_fifo_deq;
  wire [16-1:0] _mul_15_x_source_fifo_rdata;
  reg [16-1:0] _mul_15_x_source_empty_data;
  reg _mul_15_y_idle;
  reg [33-1:0] _mul_15_y_source_count;
  reg [5-1:0] _mul_15_y_source_mode;
  reg [16-1:0] _mul_15_y_source_generator_id;
  reg [32-1:0] _mul_15_y_source_offset;
  reg [33-1:0] _mul_15_y_source_size;
  reg [32-1:0] _mul_15_y_source_stride;
  reg [32-1:0] _mul_15_y_source_offset_buf;
  reg [33-1:0] _mul_15_y_source_size_buf;
  reg [32-1:0] _mul_15_y_source_stride_buf;
  reg [8-1:0] _mul_15_y_source_sel;
  reg [32-1:0] _mul_15_y_source_ram_raddr;
  reg _mul_15_y_source_ram_renable;
  wire [16-1:0] _mul_15_y_source_ram_rdata;
  reg _mul_15_y_source_fifo_deq;
  wire [16-1:0] _mul_15_y_source_fifo_rdata;
  reg [16-1:0] _mul_15_y_source_empty_data;
  reg _mul_15_rshift_idle;
  reg [33-1:0] _mul_15_rshift_source_count;
  reg [5-1:0] _mul_15_rshift_source_mode;
  reg [16-1:0] _mul_15_rshift_source_generator_id;
  reg [32-1:0] _mul_15_rshift_source_offset;
  reg [33-1:0] _mul_15_rshift_source_size;
  reg [32-1:0] _mul_15_rshift_source_stride;
  reg [32-1:0] _mul_15_rshift_source_offset_buf;
  reg [33-1:0] _mul_15_rshift_source_size_buf;
  reg [32-1:0] _mul_15_rshift_source_stride_buf;
  reg [8-1:0] _mul_15_rshift_source_sel;
  reg [32-1:0] _mul_15_rshift_source_ram_raddr;
  reg _mul_15_rshift_source_ram_renable;
  wire [32-1:0] _mul_15_rshift_source_ram_rdata;
  reg _mul_15_rshift_source_fifo_deq;
  wire [32-1:0] _mul_15_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_15_rshift_source_empty_data;
  reg [33-1:0] _mul_15_z_sink_count;
  reg [5-1:0] _mul_15_z_sink_mode;
  reg [16-1:0] _mul_15_z_sink_generator_id;
  reg [32-1:0] _mul_15_z_sink_offset;
  reg [33-1:0] _mul_15_z_sink_size;
  reg [32-1:0] _mul_15_z_sink_stride;
  reg [32-1:0] _mul_15_z_sink_offset_buf;
  reg [33-1:0] _mul_15_z_sink_size_buf;
  reg [32-1:0] _mul_15_z_sink_stride_buf;
  reg [8-1:0] _mul_15_z_sink_sel;
  reg [32-1:0] _mul_15_z_sink_waddr;
  reg _mul_15_z_sink_wenable;
  reg [32-1:0] _mul_15_z_sink_wdata;
  reg _mul_15_z_sink_fifo_enq;
  reg [32-1:0] _mul_15_z_sink_fifo_wdata;
  reg [32-1:0] _mul_15_z_sink_immediate;
  reg _mul_16_stream_ivalid;
  wire _mul_16_stream_oready;
  wire _mul_16_stream_internal_oready;
  assign _mul_16_stream_internal_oready = 1;
  reg [32-1:0] _mul_16_fsm;
  localparam _mul_16_fsm_init = 0;
  wire _mul_16_run_flag;
  assign _mul_16_run_flag = 0;
  reg _mul_16_source_start;
  wire _mul_16_source_stop;
  reg _mul_16_source_busy;
  wire _mul_16_sink_start;
  wire _mul_16_sink_stop;
  wire _mul_16_sink_busy;
  wire _mul_16_busy;
  reg _mul_16_busy_reg;
  wire _mul_16_is_root;
  reg _mul_16_x_idle;
  reg [33-1:0] _mul_16_x_source_count;
  reg [5-1:0] _mul_16_x_source_mode;
  reg [16-1:0] _mul_16_x_source_generator_id;
  reg [32-1:0] _mul_16_x_source_offset;
  reg [33-1:0] _mul_16_x_source_size;
  reg [32-1:0] _mul_16_x_source_stride;
  reg [32-1:0] _mul_16_x_source_offset_buf;
  reg [33-1:0] _mul_16_x_source_size_buf;
  reg [32-1:0] _mul_16_x_source_stride_buf;
  reg [8-1:0] _mul_16_x_source_sel;
  reg [32-1:0] _mul_16_x_source_ram_raddr;
  reg _mul_16_x_source_ram_renable;
  wire [16-1:0] _mul_16_x_source_ram_rdata;
  reg _mul_16_x_source_fifo_deq;
  wire [16-1:0] _mul_16_x_source_fifo_rdata;
  reg [16-1:0] _mul_16_x_source_empty_data;
  reg _mul_16_y_idle;
  reg [33-1:0] _mul_16_y_source_count;
  reg [5-1:0] _mul_16_y_source_mode;
  reg [16-1:0] _mul_16_y_source_generator_id;
  reg [32-1:0] _mul_16_y_source_offset;
  reg [33-1:0] _mul_16_y_source_size;
  reg [32-1:0] _mul_16_y_source_stride;
  reg [32-1:0] _mul_16_y_source_offset_buf;
  reg [33-1:0] _mul_16_y_source_size_buf;
  reg [32-1:0] _mul_16_y_source_stride_buf;
  reg [8-1:0] _mul_16_y_source_sel;
  reg [32-1:0] _mul_16_y_source_ram_raddr;
  reg _mul_16_y_source_ram_renable;
  wire [16-1:0] _mul_16_y_source_ram_rdata;
  reg _mul_16_y_source_fifo_deq;
  wire [16-1:0] _mul_16_y_source_fifo_rdata;
  reg [16-1:0] _mul_16_y_source_empty_data;
  reg _mul_16_rshift_idle;
  reg [33-1:0] _mul_16_rshift_source_count;
  reg [5-1:0] _mul_16_rshift_source_mode;
  reg [16-1:0] _mul_16_rshift_source_generator_id;
  reg [32-1:0] _mul_16_rshift_source_offset;
  reg [33-1:0] _mul_16_rshift_source_size;
  reg [32-1:0] _mul_16_rshift_source_stride;
  reg [32-1:0] _mul_16_rshift_source_offset_buf;
  reg [33-1:0] _mul_16_rshift_source_size_buf;
  reg [32-1:0] _mul_16_rshift_source_stride_buf;
  reg [8-1:0] _mul_16_rshift_source_sel;
  reg [32-1:0] _mul_16_rshift_source_ram_raddr;
  reg _mul_16_rshift_source_ram_renable;
  wire [32-1:0] _mul_16_rshift_source_ram_rdata;
  reg _mul_16_rshift_source_fifo_deq;
  wire [32-1:0] _mul_16_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_16_rshift_source_empty_data;
  reg [33-1:0] _mul_16_z_sink_count;
  reg [5-1:0] _mul_16_z_sink_mode;
  reg [16-1:0] _mul_16_z_sink_generator_id;
  reg [32-1:0] _mul_16_z_sink_offset;
  reg [33-1:0] _mul_16_z_sink_size;
  reg [32-1:0] _mul_16_z_sink_stride;
  reg [32-1:0] _mul_16_z_sink_offset_buf;
  reg [33-1:0] _mul_16_z_sink_size_buf;
  reg [32-1:0] _mul_16_z_sink_stride_buf;
  reg [8-1:0] _mul_16_z_sink_sel;
  reg [32-1:0] _mul_16_z_sink_waddr;
  reg _mul_16_z_sink_wenable;
  reg [32-1:0] _mul_16_z_sink_wdata;
  reg _mul_16_z_sink_fifo_enq;
  reg [32-1:0] _mul_16_z_sink_fifo_wdata;
  reg [32-1:0] _mul_16_z_sink_immediate;
  reg __reduce_max_17_stream_ivalid;
  wire __reduce_max_17_stream_oready;
  wire __reduce_max_17_stream_internal_oready;
  assign __reduce_max_17_stream_internal_oready = 1;
  reg [32-1:0] __reduce_max_17_fsm;
  localparam __reduce_max_17_fsm_init = 0;
  wire __reduce_max_17_run_flag;
  assign __reduce_max_17_run_flag = 0;
  reg __reduce_max_17_source_start;
  wire __reduce_max_17_source_stop;
  reg __reduce_max_17_source_busy;
  wire __reduce_max_17_sink_start;
  wire __reduce_max_17_sink_stop;
  wire __reduce_max_17_sink_busy;
  wire __reduce_max_17_busy;
  reg __reduce_max_17_busy_reg;
  wire __reduce_max_17_is_root;
  reg __reduce_max_17_x_idle;
  reg [33-1:0] __reduce_max_17_x_source_count;
  reg [5-1:0] __reduce_max_17_x_source_mode;
  reg [16-1:0] __reduce_max_17_x_source_generator_id;
  reg [32-1:0] __reduce_max_17_x_source_offset;
  reg [33-1:0] __reduce_max_17_x_source_size;
  reg [32-1:0] __reduce_max_17_x_source_stride;
  reg [32-1:0] __reduce_max_17_x_source_offset_buf;
  reg [33-1:0] __reduce_max_17_x_source_size_buf;
  reg [32-1:0] __reduce_max_17_x_source_stride_buf;
  reg [8-1:0] __reduce_max_17_x_source_sel;
  reg [32-1:0] __reduce_max_17_x_source_ram_raddr;
  reg __reduce_max_17_x_source_ram_renable;
  wire [16-1:0] __reduce_max_17_x_source_ram_rdata;
  reg __reduce_max_17_x_source_fifo_deq;
  wire [16-1:0] __reduce_max_17_x_source_fifo_rdata;
  reg [16-1:0] __reduce_max_17_x_source_empty_data;
  reg [32-1:0] __reduce_max_17_size_next_parameter_data;
  reg [33-1:0] __reduce_max_17_data_sink_count;
  reg [5-1:0] __reduce_max_17_data_sink_mode;
  reg [16-1:0] __reduce_max_17_data_sink_generator_id;
  reg [32-1:0] __reduce_max_17_data_sink_offset;
  reg [33-1:0] __reduce_max_17_data_sink_size;
  reg [32-1:0] __reduce_max_17_data_sink_stride;
  reg [32-1:0] __reduce_max_17_data_sink_offset_buf;
  reg [33-1:0] __reduce_max_17_data_sink_size_buf;
  reg [32-1:0] __reduce_max_17_data_sink_stride_buf;
  reg [8-1:0] __reduce_max_17_data_sink_sel;
  reg [32-1:0] __reduce_max_17_data_sink_waddr;
  reg __reduce_max_17_data_sink_wenable;
  reg [16-1:0] __reduce_max_17_data_sink_wdata;
  reg __reduce_max_17_data_sink_fifo_enq;
  reg [16-1:0] __reduce_max_17_data_sink_fifo_wdata;
  reg [16-1:0] __reduce_max_17_data_sink_immediate;
  reg [33-1:0] __reduce_max_17_valid_sink_count;
  reg [5-1:0] __reduce_max_17_valid_sink_mode;
  reg [16-1:0] __reduce_max_17_valid_sink_generator_id;
  reg [32-1:0] __reduce_max_17_valid_sink_offset;
  reg [33-1:0] __reduce_max_17_valid_sink_size;
  reg [32-1:0] __reduce_max_17_valid_sink_stride;
  reg [32-1:0] __reduce_max_17_valid_sink_offset_buf;
  reg [33-1:0] __reduce_max_17_valid_sink_size_buf;
  reg [32-1:0] __reduce_max_17_valid_sink_stride_buf;
  reg [8-1:0] __reduce_max_17_valid_sink_sel;
  reg [32-1:0] __reduce_max_17_valid_sink_waddr;
  reg __reduce_max_17_valid_sink_wenable;
  reg [1-1:0] __reduce_max_17_valid_sink_wdata;
  reg __reduce_max_17_valid_sink_fifo_enq;
  reg [1-1:0] __reduce_max_17_valid_sink_fifo_wdata;
  reg [1-1:0] __reduce_max_17_valid_sink_immediate;
  reg __reduce_max_18_stream_ivalid;
  wire __reduce_max_18_stream_oready;
  wire __reduce_max_18_stream_internal_oready;
  assign __reduce_max_18_stream_internal_oready = 1;
  reg [32-1:0] __reduce_max_18_fsm;
  localparam __reduce_max_18_fsm_init = 0;
  wire __reduce_max_18_run_flag;
  assign __reduce_max_18_run_flag = 0;
  reg __reduce_max_18_source_start;
  wire __reduce_max_18_source_stop;
  reg __reduce_max_18_source_busy;
  wire __reduce_max_18_sink_start;
  wire __reduce_max_18_sink_stop;
  wire __reduce_max_18_sink_busy;
  wire __reduce_max_18_busy;
  reg __reduce_max_18_busy_reg;
  wire __reduce_max_18_is_root;
  reg __reduce_max_18_x_idle;
  reg [33-1:0] __reduce_max_18_x_source_count;
  reg [5-1:0] __reduce_max_18_x_source_mode;
  reg [16-1:0] __reduce_max_18_x_source_generator_id;
  reg [32-1:0] __reduce_max_18_x_source_offset;
  reg [33-1:0] __reduce_max_18_x_source_size;
  reg [32-1:0] __reduce_max_18_x_source_stride;
  reg [32-1:0] __reduce_max_18_x_source_offset_buf;
  reg [33-1:0] __reduce_max_18_x_source_size_buf;
  reg [32-1:0] __reduce_max_18_x_source_stride_buf;
  reg [8-1:0] __reduce_max_18_x_source_sel;
  reg [32-1:0] __reduce_max_18_x_source_ram_raddr;
  reg __reduce_max_18_x_source_ram_renable;
  wire [16-1:0] __reduce_max_18_x_source_ram_rdata;
  reg __reduce_max_18_x_source_fifo_deq;
  wire [16-1:0] __reduce_max_18_x_source_fifo_rdata;
  reg [16-1:0] __reduce_max_18_x_source_empty_data;
  reg [32-1:0] __reduce_max_18_size_next_parameter_data;
  reg [33-1:0] __reduce_max_18_data_sink_count;
  reg [5-1:0] __reduce_max_18_data_sink_mode;
  reg [16-1:0] __reduce_max_18_data_sink_generator_id;
  reg [32-1:0] __reduce_max_18_data_sink_offset;
  reg [33-1:0] __reduce_max_18_data_sink_size;
  reg [32-1:0] __reduce_max_18_data_sink_stride;
  reg [32-1:0] __reduce_max_18_data_sink_offset_buf;
  reg [33-1:0] __reduce_max_18_data_sink_size_buf;
  reg [32-1:0] __reduce_max_18_data_sink_stride_buf;
  reg [8-1:0] __reduce_max_18_data_sink_sel;
  reg [32-1:0] __reduce_max_18_data_sink_waddr;
  reg __reduce_max_18_data_sink_wenable;
  reg [16-1:0] __reduce_max_18_data_sink_wdata;
  reg __reduce_max_18_data_sink_fifo_enq;
  reg [16-1:0] __reduce_max_18_data_sink_fifo_wdata;
  reg [16-1:0] __reduce_max_18_data_sink_immediate;
  reg [33-1:0] __reduce_max_18_valid_sink_count;
  reg [5-1:0] __reduce_max_18_valid_sink_mode;
  reg [16-1:0] __reduce_max_18_valid_sink_generator_id;
  reg [32-1:0] __reduce_max_18_valid_sink_offset;
  reg [33-1:0] __reduce_max_18_valid_sink_size;
  reg [32-1:0] __reduce_max_18_valid_sink_stride;
  reg [32-1:0] __reduce_max_18_valid_sink_offset_buf;
  reg [33-1:0] __reduce_max_18_valid_sink_size_buf;
  reg [32-1:0] __reduce_max_18_valid_sink_stride_buf;
  reg [8-1:0] __reduce_max_18_valid_sink_sel;
  reg [32-1:0] __reduce_max_18_valid_sink_waddr;
  reg __reduce_max_18_valid_sink_wenable;
  reg [1-1:0] __reduce_max_18_valid_sink_wdata;
  reg __reduce_max_18_valid_sink_fifo_enq;
  reg [1-1:0] __reduce_max_18_valid_sink_fifo_wdata;
  reg [1-1:0] __reduce_max_18_valid_sink_immediate;
  reg _stream_conv2d_4_stream_ivalid;
  wire _stream_conv2d_4_stream_oready;
  wire _stream_conv2d_4_stream_internal_oready;
  assign _stream_conv2d_4_stream_oready = _stream_conv2d_4_stream_internal_oready;
  reg [32-1:0] _stream_conv2d_4_fsm;
  localparam _stream_conv2d_4_fsm_init = 0;
  wire _stream_conv2d_4_run_flag;
  reg _stream_conv2d_4_source_start;
  wire _stream_conv2d_4_source_stop;
  reg _stream_conv2d_4_source_busy;
  wire _stream_conv2d_4_sink_start;
  wire _stream_conv2d_4_sink_stop;
  wire _stream_conv2d_4_sink_busy;
  wire _stream_conv2d_4_busy;
  reg _stream_conv2d_4_busy_reg;
  wire _stream_conv2d_4_is_root;
  assign _stream_conv2d_4_is_root = 1;
  reg [8-1:0] _stream_conv2d_4_parameter_0_next_parameter_data;
  reg [2-1:0] _stream_conv2d_4_parameter_1_next_parameter_data;
  reg [2-1:0] _stream_conv2d_4_parameter_2_next_parameter_data;
  reg [9-1:0] _stream_conv2d_4_parameter_3_next_parameter_data;
  reg [1-1:0] _stream_conv2d_4_parameter_4_next_parameter_data;
  reg [1-1:0] _stream_conv2d_4_parameter_6_next_parameter_data;
  reg _stream_conv2d_4_source_7_idle;
  reg [33-1:0] _stream_conv2d_4_source_7_source_count;
  reg [5-1:0] _stream_conv2d_4_source_7_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_7_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_7_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_7_source_size;
  reg [32-1:0] _stream_conv2d_4_source_7_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_7_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_7_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_7_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_7_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_7_source_ram_raddr;
  reg _stream_conv2d_4_source_7_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_7_source_ram_rdata;
  reg _stream_conv2d_4_source_7_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_7_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_7_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_8_next_parameter_data;
  reg _stream_conv2d_4_source_9_idle;
  reg [33-1:0] _stream_conv2d_4_source_9_source_count;
  reg [5-1:0] _stream_conv2d_4_source_9_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_9_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_9_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_9_source_size;
  reg [32-1:0] _stream_conv2d_4_source_9_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_9_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_9_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_9_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_9_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_9_source_ram_raddr;
  reg _stream_conv2d_4_source_9_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_9_source_ram_rdata;
  reg _stream_conv2d_4_source_9_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_9_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_9_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_10_next_parameter_data;
  reg _stream_conv2d_4_source_11_idle;
  reg [33-1:0] _stream_conv2d_4_source_11_source_count;
  reg [5-1:0] _stream_conv2d_4_source_11_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_11_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_11_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_11_source_size;
  reg [32-1:0] _stream_conv2d_4_source_11_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_11_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_11_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_11_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_11_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_11_source_ram_raddr;
  reg _stream_conv2d_4_source_11_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_11_source_ram_rdata;
  reg _stream_conv2d_4_source_11_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_11_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_11_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_12_next_parameter_data;
  reg _stream_conv2d_4_source_13_idle;
  reg [33-1:0] _stream_conv2d_4_source_13_source_count;
  reg [5-1:0] _stream_conv2d_4_source_13_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_13_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_13_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_13_source_size;
  reg [32-1:0] _stream_conv2d_4_source_13_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_13_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_13_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_13_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_13_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_13_source_ram_raddr;
  reg _stream_conv2d_4_source_13_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_13_source_ram_rdata;
  reg _stream_conv2d_4_source_13_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_13_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_13_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_14_next_parameter_data;
  reg _stream_conv2d_4_source_15_idle;
  reg [33-1:0] _stream_conv2d_4_source_15_source_count;
  reg [5-1:0] _stream_conv2d_4_source_15_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_15_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_15_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_15_source_size;
  reg [32-1:0] _stream_conv2d_4_source_15_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_15_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_15_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_15_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_15_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_15_source_ram_raddr;
  reg _stream_conv2d_4_source_15_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_15_source_ram_rdata;
  reg _stream_conv2d_4_source_15_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_15_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_15_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_16_next_parameter_data;
  reg [1-1:0] _stream_conv2d_4_parameter_17_next_parameter_data;
  reg [1-1:0] _stream_conv2d_4_parameter_18_next_parameter_data;
  reg [1-1:0] _stream_conv2d_4_parameter_19_next_parameter_data;
  reg _stream_conv2d_4_source_20_idle;
  reg [33-1:0] _stream_conv2d_4_source_20_source_count;
  reg [5-1:0] _stream_conv2d_4_source_20_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_20_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_20_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_20_source_size;
  reg [32-1:0] _stream_conv2d_4_source_20_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_20_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_20_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_20_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_20_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_20_source_ram_raddr;
  reg _stream_conv2d_4_source_20_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_20_source_ram_rdata;
  reg _stream_conv2d_4_source_20_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_20_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_20_source_empty_data;
  reg _stream_conv2d_4_source_21_idle;
  reg [33-1:0] _stream_conv2d_4_source_21_source_count;
  reg [5-1:0] _stream_conv2d_4_source_21_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_21_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_21_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_21_source_size;
  reg [32-1:0] _stream_conv2d_4_source_21_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_21_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_21_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_21_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_21_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_21_source_ram_raddr;
  reg _stream_conv2d_4_source_21_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_21_source_ram_rdata;
  reg _stream_conv2d_4_source_21_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_21_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_21_source_empty_data;
  reg _stream_conv2d_4_source_22_idle;
  reg [33-1:0] _stream_conv2d_4_source_22_source_count;
  reg [5-1:0] _stream_conv2d_4_source_22_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_22_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_22_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_22_source_size;
  reg [32-1:0] _stream_conv2d_4_source_22_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_22_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_22_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_22_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_22_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_22_source_ram_raddr;
  reg _stream_conv2d_4_source_22_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_22_source_ram_rdata;
  reg _stream_conv2d_4_source_22_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_22_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_22_source_empty_data;
  reg _stream_conv2d_4_source_23_idle;
  reg [33-1:0] _stream_conv2d_4_source_23_source_count;
  reg [5-1:0] _stream_conv2d_4_source_23_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_23_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_23_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_23_source_size;
  reg [32-1:0] _stream_conv2d_4_source_23_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_23_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_23_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_23_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_23_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_23_source_ram_raddr;
  reg _stream_conv2d_4_source_23_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_23_source_ram_rdata;
  reg _stream_conv2d_4_source_23_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_23_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_23_source_empty_data;
  reg _stream_conv2d_4_source_24_idle;
  reg [33-1:0] _stream_conv2d_4_source_24_source_count;
  reg [5-1:0] _stream_conv2d_4_source_24_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_24_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_24_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_24_source_size;
  reg [32-1:0] _stream_conv2d_4_source_24_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_24_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_24_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_24_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_24_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_24_source_ram_raddr;
  reg _stream_conv2d_4_source_24_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_24_source_ram_rdata;
  reg _stream_conv2d_4_source_24_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_24_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_24_source_empty_data;
  reg _stream_conv2d_4_source_25_idle;
  reg [33-1:0] _stream_conv2d_4_source_25_source_count;
  reg [5-1:0] _stream_conv2d_4_source_25_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_25_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_25_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_25_source_size;
  reg [32-1:0] _stream_conv2d_4_source_25_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_25_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_25_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_25_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_25_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_25_source_ram_raddr;
  reg _stream_conv2d_4_source_25_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_25_source_ram_rdata;
  reg _stream_conv2d_4_source_25_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_25_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_25_source_empty_data;
  reg _stream_conv2d_4_source_26_idle;
  reg [33-1:0] _stream_conv2d_4_source_26_source_count;
  reg [5-1:0] _stream_conv2d_4_source_26_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_26_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_26_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_26_source_size;
  reg [32-1:0] _stream_conv2d_4_source_26_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_26_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_26_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_26_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_26_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_26_source_ram_raddr;
  reg _stream_conv2d_4_source_26_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_26_source_ram_rdata;
  reg _stream_conv2d_4_source_26_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_26_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_26_source_empty_data;
  reg _stream_conv2d_4_source_27_idle;
  reg [33-1:0] _stream_conv2d_4_source_27_source_count;
  reg [5-1:0] _stream_conv2d_4_source_27_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_27_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_27_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_27_source_size;
  reg [32-1:0] _stream_conv2d_4_source_27_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_27_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_27_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_27_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_27_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_27_source_ram_raddr;
  reg _stream_conv2d_4_source_27_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_27_source_ram_rdata;
  reg _stream_conv2d_4_source_27_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_27_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_27_source_empty_data;
  reg _stream_conv2d_4_source_28_idle;
  reg [33-1:0] _stream_conv2d_4_source_28_source_count;
  reg [5-1:0] _stream_conv2d_4_source_28_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_28_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_28_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_28_source_size;
  reg [32-1:0] _stream_conv2d_4_source_28_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_28_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_28_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_28_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_28_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_28_source_ram_raddr;
  reg _stream_conv2d_4_source_28_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_28_source_ram_rdata;
  reg _stream_conv2d_4_source_28_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_28_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_28_source_empty_data;
  reg _stream_conv2d_4_source_29_idle;
  reg [33-1:0] _stream_conv2d_4_source_29_source_count;
  reg [5-1:0] _stream_conv2d_4_source_29_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_29_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_29_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_29_source_size;
  reg [32-1:0] _stream_conv2d_4_source_29_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_29_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_29_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_29_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_29_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_29_source_ram_raddr;
  reg _stream_conv2d_4_source_29_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_29_source_ram_rdata;
  reg _stream_conv2d_4_source_29_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_29_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_29_source_empty_data;
  reg _stream_conv2d_4_source_30_idle;
  reg [33-1:0] _stream_conv2d_4_source_30_source_count;
  reg [5-1:0] _stream_conv2d_4_source_30_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_30_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_30_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_30_source_size;
  reg [32-1:0] _stream_conv2d_4_source_30_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_30_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_30_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_30_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_30_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_30_source_ram_raddr;
  reg _stream_conv2d_4_source_30_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_30_source_ram_rdata;
  reg _stream_conv2d_4_source_30_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_30_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_30_source_empty_data;
  reg _stream_conv2d_4_source_31_idle;
  reg [33-1:0] _stream_conv2d_4_source_31_source_count;
  reg [5-1:0] _stream_conv2d_4_source_31_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_31_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_31_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_31_source_size;
  reg [32-1:0] _stream_conv2d_4_source_31_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_31_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_31_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_31_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_31_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_31_source_ram_raddr;
  reg _stream_conv2d_4_source_31_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_31_source_ram_rdata;
  reg _stream_conv2d_4_source_31_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_31_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_31_source_empty_data;
  reg _stream_conv2d_4_source_32_idle;
  reg [33-1:0] _stream_conv2d_4_source_32_source_count;
  reg [5-1:0] _stream_conv2d_4_source_32_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_32_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_32_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_32_source_size;
  reg [32-1:0] _stream_conv2d_4_source_32_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_32_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_32_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_32_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_32_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_32_source_ram_raddr;
  reg _stream_conv2d_4_source_32_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_32_source_ram_rdata;
  reg _stream_conv2d_4_source_32_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_32_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_32_source_empty_data;
  reg _stream_conv2d_4_source_33_idle;
  reg [33-1:0] _stream_conv2d_4_source_33_source_count;
  reg [5-1:0] _stream_conv2d_4_source_33_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_33_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_33_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_33_source_size;
  reg [32-1:0] _stream_conv2d_4_source_33_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_33_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_33_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_33_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_33_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_33_source_ram_raddr;
  reg _stream_conv2d_4_source_33_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_33_source_ram_rdata;
  reg _stream_conv2d_4_source_33_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_33_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_33_source_empty_data;
  reg _stream_conv2d_4_source_34_idle;
  reg [33-1:0] _stream_conv2d_4_source_34_source_count;
  reg [5-1:0] _stream_conv2d_4_source_34_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_34_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_34_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_34_source_size;
  reg [32-1:0] _stream_conv2d_4_source_34_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_34_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_34_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_34_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_34_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_34_source_ram_raddr;
  reg _stream_conv2d_4_source_34_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_34_source_ram_rdata;
  reg _stream_conv2d_4_source_34_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_34_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_34_source_empty_data;
  reg _stream_conv2d_4_source_35_idle;
  reg [33-1:0] _stream_conv2d_4_source_35_source_count;
  reg [5-1:0] _stream_conv2d_4_source_35_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_35_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_35_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_35_source_size;
  reg [32-1:0] _stream_conv2d_4_source_35_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_35_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_35_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_35_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_35_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_35_source_ram_raddr;
  reg _stream_conv2d_4_source_35_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_35_source_ram_rdata;
  reg _stream_conv2d_4_source_35_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_35_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_35_source_empty_data;
  reg _stream_conv2d_4_source_36_idle;
  reg [33-1:0] _stream_conv2d_4_source_36_source_count;
  reg [5-1:0] _stream_conv2d_4_source_36_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_36_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_36_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_36_source_size;
  reg [32-1:0] _stream_conv2d_4_source_36_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_36_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_36_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_36_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_36_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_36_source_ram_raddr;
  reg _stream_conv2d_4_source_36_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_36_source_ram_rdata;
  reg _stream_conv2d_4_source_36_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_36_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_36_source_empty_data;
  reg _stream_conv2d_4_source_37_idle;
  reg [33-1:0] _stream_conv2d_4_source_37_source_count;
  reg [5-1:0] _stream_conv2d_4_source_37_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_37_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_37_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_37_source_size;
  reg [32-1:0] _stream_conv2d_4_source_37_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_37_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_37_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_37_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_37_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_37_source_ram_raddr;
  reg _stream_conv2d_4_source_37_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_37_source_ram_rdata;
  reg _stream_conv2d_4_source_37_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_37_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_37_source_empty_data;
  wire signed [16-1:0] mul_8_x_data;
  wire signed [16-1:0] mul_8_y_data;
  wire [5-1:0] mul_8_rshift_data;
  reg __mul_8_stream_ivalid_1;
  reg __mul_8_stream_ivalid_2;
  reg __mul_8_stream_ivalid_3;
  reg __mul_8_stream_ivalid_4;
  reg __mul_8_stream_ivalid_5;
  reg __mul_8_stream_ivalid_6;
  reg __mul_8_stream_ivalid_7;
  reg __mul_8_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_139;
  reg [5-1:0] _minus_data_141;
  reg [1-1:0] _greatereq_data_152;
  reg signed [16-1:0] __delay_data_721__variable_136;
  reg signed [16-1:0] __delay_data_724__variable_137;
  reg [5-1:0] __delay_data_727__variable_138;
  reg signed [34-1:0] _sll_data_143;
  reg [1-1:0] __delay_data_718_greaterthan_139;
  reg [1-1:0] __delay_data_719_greatereq_152;
  reg signed [16-1:0] __delay_data_722__delay_721__variable_136;
  reg signed [16-1:0] __delay_data_725__delay_724__variable_137;
  reg [5-1:0] __delay_data_728__delay_727__variable_138;
  reg signed [32-1:0] _cond_data_149;
  reg [1-1:0] __delay_data_720__delay_719_greatereq_152;
  reg signed [16-1:0] __delay_data_723__delay_722__delay_721__variable_136;
  reg signed [16-1:0] __delay_data_726__delay_725__delay_724__variable_137;
  reg [5-1:0] __delay_data_729__delay_728__delay_727__variable_138;
  wire signed [16-1:0] _uminus_data_151;
  assign _uminus_data_151 = -_cond_data_149;
  wire signed [16-1:0] _cond_data_154;
  assign _cond_data_154 = (__delay_data_720__delay_719_greatereq_152)? _cond_data_149 : _uminus_data_151;
  wire signed [32-1:0] __muladd_madd_odata_155;
  reg signed [32-1:0] __muladd_madd_odata_reg_155;
  wire signed [32-1:0] __muladd_data_155;
  assign __muladd_data_155 = __muladd_madd_odata_reg_155;
  wire __muladd_madd_update_155;
  assign __muladd_madd_update_155 = _mul_8_stream_oready;

  madd_0
  __muladd_madd_155
  (
    .CLK(CLK),
    .update(__muladd_madd_update_155),
    .a(__delay_data_723__delay_722__delay_721__variable_136),
    .b(__delay_data_726__delay_725__delay_724__variable_137),
    .c(_cond_data_154),
    .d(__muladd_madd_odata_155)
  );

  reg [5-1:0] __delay_data_730__delay_729__delay_728____variable_138;
  reg [5-1:0] __delay_data_731__delay_730__delay_729____variable_138;
  reg [5-1:0] __delay_data_732__delay_731__delay_730____variable_138;
  reg [5-1:0] __delay_data_733__delay_732__delay_731____variable_138;
  reg signed [32-1:0] _sra_data_156;
  wire signed [32-1:0] mul_8_z_data;
  assign mul_8_z_data = _sra_data_156;
  wire signed [16-1:0] mul_9_x_data;
  wire signed [16-1:0] mul_9_y_data;
  wire [5-1:0] mul_9_rshift_data;
  reg __mul_9_stream_ivalid_1;
  reg __mul_9_stream_ivalid_2;
  reg __mul_9_stream_ivalid_3;
  reg __mul_9_stream_ivalid_4;
  reg __mul_9_stream_ivalid_5;
  reg __mul_9_stream_ivalid_6;
  reg __mul_9_stream_ivalid_7;
  reg __mul_9_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_160;
  reg [5-1:0] _minus_data_162;
  reg [1-1:0] _greatereq_data_173;
  reg signed [16-1:0] __delay_data_740__variable_157;
  reg signed [16-1:0] __delay_data_743__variable_158;
  reg [5-1:0] __delay_data_746__variable_159;
  reg signed [34-1:0] _sll_data_164;
  reg [1-1:0] __delay_data_737_greaterthan_160;
  reg [1-1:0] __delay_data_738_greatereq_173;
  reg signed [16-1:0] __delay_data_741__delay_740__variable_157;
  reg signed [16-1:0] __delay_data_744__delay_743__variable_158;
  reg [5-1:0] __delay_data_747__delay_746__variable_159;
  reg signed [32-1:0] _cond_data_170;
  reg [1-1:0] __delay_data_739__delay_738_greatereq_173;
  reg signed [16-1:0] __delay_data_742__delay_741__delay_740__variable_157;
  reg signed [16-1:0] __delay_data_745__delay_744__delay_743__variable_158;
  reg [5-1:0] __delay_data_748__delay_747__delay_746__variable_159;
  wire signed [16-1:0] _uminus_data_172;
  assign _uminus_data_172 = -_cond_data_170;
  wire signed [16-1:0] _cond_data_175;
  assign _cond_data_175 = (__delay_data_739__delay_738_greatereq_173)? _cond_data_170 : _uminus_data_172;
  wire signed [32-1:0] __muladd_madd_odata_176;
  reg signed [32-1:0] __muladd_madd_odata_reg_176;
  wire signed [32-1:0] __muladd_data_176;
  assign __muladd_data_176 = __muladd_madd_odata_reg_176;
  wire __muladd_madd_update_176;
  assign __muladd_madd_update_176 = _mul_9_stream_oready;

  madd_1
  __muladd_madd_176
  (
    .CLK(CLK),
    .update(__muladd_madd_update_176),
    .a(__delay_data_742__delay_741__delay_740__variable_157),
    .b(__delay_data_745__delay_744__delay_743__variable_158),
    .c(_cond_data_175),
    .d(__muladd_madd_odata_176)
  );

  reg [5-1:0] __delay_data_749__delay_748__delay_747____variable_159;
  reg [5-1:0] __delay_data_750__delay_749__delay_748____variable_159;
  reg [5-1:0] __delay_data_751__delay_750__delay_749____variable_159;
  reg [5-1:0] __delay_data_752__delay_751__delay_750____variable_159;
  reg signed [32-1:0] _sra_data_177;
  wire signed [32-1:0] mul_9_z_data;
  assign mul_9_z_data = _sra_data_177;
  wire signed [16-1:0] mul_10_x_data;
  wire signed [16-1:0] mul_10_y_data;
  wire [5-1:0] mul_10_rshift_data;
  reg __mul_10_stream_ivalid_1;
  reg __mul_10_stream_ivalid_2;
  reg __mul_10_stream_ivalid_3;
  reg __mul_10_stream_ivalid_4;
  reg __mul_10_stream_ivalid_5;
  reg __mul_10_stream_ivalid_6;
  reg __mul_10_stream_ivalid_7;
  reg __mul_10_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_181;
  reg [5-1:0] _minus_data_183;
  reg [1-1:0] _greatereq_data_194;
  reg signed [16-1:0] __delay_data_759__variable_178;
  reg signed [16-1:0] __delay_data_762__variable_179;
  reg [5-1:0] __delay_data_765__variable_180;
  reg signed [34-1:0] _sll_data_185;
  reg [1-1:0] __delay_data_756_greaterthan_181;
  reg [1-1:0] __delay_data_757_greatereq_194;
  reg signed [16-1:0] __delay_data_760__delay_759__variable_178;
  reg signed [16-1:0] __delay_data_763__delay_762__variable_179;
  reg [5-1:0] __delay_data_766__delay_765__variable_180;
  reg signed [32-1:0] _cond_data_191;
  reg [1-1:0] __delay_data_758__delay_757_greatereq_194;
  reg signed [16-1:0] __delay_data_761__delay_760__delay_759__variable_178;
  reg signed [16-1:0] __delay_data_764__delay_763__delay_762__variable_179;
  reg [5-1:0] __delay_data_767__delay_766__delay_765__variable_180;
  wire signed [16-1:0] _uminus_data_193;
  assign _uminus_data_193 = -_cond_data_191;
  wire signed [16-1:0] _cond_data_196;
  assign _cond_data_196 = (__delay_data_758__delay_757_greatereq_194)? _cond_data_191 : _uminus_data_193;
  wire signed [32-1:0] __muladd_madd_odata_197;
  reg signed [32-1:0] __muladd_madd_odata_reg_197;
  wire signed [32-1:0] __muladd_data_197;
  assign __muladd_data_197 = __muladd_madd_odata_reg_197;
  wire __muladd_madd_update_197;
  assign __muladd_madd_update_197 = _mul_10_stream_oready;

  madd_2
  __muladd_madd_197
  (
    .CLK(CLK),
    .update(__muladd_madd_update_197),
    .a(__delay_data_761__delay_760__delay_759__variable_178),
    .b(__delay_data_764__delay_763__delay_762__variable_179),
    .c(_cond_data_196),
    .d(__muladd_madd_odata_197)
  );

  reg [5-1:0] __delay_data_768__delay_767__delay_766____variable_180;
  reg [5-1:0] __delay_data_769__delay_768__delay_767____variable_180;
  reg [5-1:0] __delay_data_770__delay_769__delay_768____variable_180;
  reg [5-1:0] __delay_data_771__delay_770__delay_769____variable_180;
  reg signed [32-1:0] _sra_data_198;
  wire signed [32-1:0] mul_10_z_data;
  assign mul_10_z_data = _sra_data_198;
  wire signed [16-1:0] mul_11_x_data;
  wire signed [16-1:0] mul_11_y_data;
  wire [5-1:0] mul_11_rshift_data;
  reg __mul_11_stream_ivalid_1;
  reg __mul_11_stream_ivalid_2;
  reg __mul_11_stream_ivalid_3;
  reg __mul_11_stream_ivalid_4;
  reg __mul_11_stream_ivalid_5;
  reg __mul_11_stream_ivalid_6;
  reg __mul_11_stream_ivalid_7;
  reg __mul_11_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_202;
  reg [5-1:0] _minus_data_204;
  reg [1-1:0] _greatereq_data_215;
  reg signed [16-1:0] __delay_data_778__variable_199;
  reg signed [16-1:0] __delay_data_781__variable_200;
  reg [5-1:0] __delay_data_784__variable_201;
  reg signed [34-1:0] _sll_data_206;
  reg [1-1:0] __delay_data_775_greaterthan_202;
  reg [1-1:0] __delay_data_776_greatereq_215;
  reg signed [16-1:0] __delay_data_779__delay_778__variable_199;
  reg signed [16-1:0] __delay_data_782__delay_781__variable_200;
  reg [5-1:0] __delay_data_785__delay_784__variable_201;
  reg signed [32-1:0] _cond_data_212;
  reg [1-1:0] __delay_data_777__delay_776_greatereq_215;
  reg signed [16-1:0] __delay_data_780__delay_779__delay_778__variable_199;
  reg signed [16-1:0] __delay_data_783__delay_782__delay_781__variable_200;
  reg [5-1:0] __delay_data_786__delay_785__delay_784__variable_201;
  wire signed [16-1:0] _uminus_data_214;
  assign _uminus_data_214 = -_cond_data_212;
  wire signed [16-1:0] _cond_data_217;
  assign _cond_data_217 = (__delay_data_777__delay_776_greatereq_215)? _cond_data_212 : _uminus_data_214;
  wire signed [32-1:0] __muladd_madd_odata_218;
  reg signed [32-1:0] __muladd_madd_odata_reg_218;
  wire signed [32-1:0] __muladd_data_218;
  assign __muladd_data_218 = __muladd_madd_odata_reg_218;
  wire __muladd_madd_update_218;
  assign __muladd_madd_update_218 = _mul_11_stream_oready;

  madd_3
  __muladd_madd_218
  (
    .CLK(CLK),
    .update(__muladd_madd_update_218),
    .a(__delay_data_780__delay_779__delay_778__variable_199),
    .b(__delay_data_783__delay_782__delay_781__variable_200),
    .c(_cond_data_217),
    .d(__muladd_madd_odata_218)
  );

  reg [5-1:0] __delay_data_787__delay_786__delay_785____variable_201;
  reg [5-1:0] __delay_data_788__delay_787__delay_786____variable_201;
  reg [5-1:0] __delay_data_789__delay_788__delay_787____variable_201;
  reg [5-1:0] __delay_data_790__delay_789__delay_788____variable_201;
  reg signed [32-1:0] _sra_data_219;
  wire signed [32-1:0] mul_11_z_data;
  assign mul_11_z_data = _sra_data_219;
  wire signed [16-1:0] mul_12_x_data;
  wire signed [16-1:0] mul_12_y_data;
  wire [5-1:0] mul_12_rshift_data;
  reg __mul_12_stream_ivalid_1;
  reg __mul_12_stream_ivalid_2;
  reg __mul_12_stream_ivalid_3;
  reg __mul_12_stream_ivalid_4;
  reg __mul_12_stream_ivalid_5;
  reg __mul_12_stream_ivalid_6;
  reg __mul_12_stream_ivalid_7;
  reg __mul_12_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_223;
  reg [5-1:0] _minus_data_225;
  reg [1-1:0] _greatereq_data_236;
  reg signed [16-1:0] __delay_data_797__variable_220;
  reg signed [16-1:0] __delay_data_800__variable_221;
  reg [5-1:0] __delay_data_803__variable_222;
  reg signed [34-1:0] _sll_data_227;
  reg [1-1:0] __delay_data_794_greaterthan_223;
  reg [1-1:0] __delay_data_795_greatereq_236;
  reg signed [16-1:0] __delay_data_798__delay_797__variable_220;
  reg signed [16-1:0] __delay_data_801__delay_800__variable_221;
  reg [5-1:0] __delay_data_804__delay_803__variable_222;
  reg signed [32-1:0] _cond_data_233;
  reg [1-1:0] __delay_data_796__delay_795_greatereq_236;
  reg signed [16-1:0] __delay_data_799__delay_798__delay_797__variable_220;
  reg signed [16-1:0] __delay_data_802__delay_801__delay_800__variable_221;
  reg [5-1:0] __delay_data_805__delay_804__delay_803__variable_222;
  wire signed [16-1:0] _uminus_data_235;
  assign _uminus_data_235 = -_cond_data_233;
  wire signed [16-1:0] _cond_data_238;
  assign _cond_data_238 = (__delay_data_796__delay_795_greatereq_236)? _cond_data_233 : _uminus_data_235;
  wire signed [32-1:0] __muladd_madd_odata_239;
  reg signed [32-1:0] __muladd_madd_odata_reg_239;
  wire signed [32-1:0] __muladd_data_239;
  assign __muladd_data_239 = __muladd_madd_odata_reg_239;
  wire __muladd_madd_update_239;
  assign __muladd_madd_update_239 = _mul_12_stream_oready;

  madd_4
  __muladd_madd_239
  (
    .CLK(CLK),
    .update(__muladd_madd_update_239),
    .a(__delay_data_799__delay_798__delay_797__variable_220),
    .b(__delay_data_802__delay_801__delay_800__variable_221),
    .c(_cond_data_238),
    .d(__muladd_madd_odata_239)
  );

  reg [5-1:0] __delay_data_806__delay_805__delay_804____variable_222;
  reg [5-1:0] __delay_data_807__delay_806__delay_805____variable_222;
  reg [5-1:0] __delay_data_808__delay_807__delay_806____variable_222;
  reg [5-1:0] __delay_data_809__delay_808__delay_807____variable_222;
  reg signed [32-1:0] _sra_data_240;
  wire signed [32-1:0] mul_12_z_data;
  assign mul_12_z_data = _sra_data_240;
  wire signed [16-1:0] mul_13_x_data;
  wire signed [16-1:0] mul_13_y_data;
  wire [5-1:0] mul_13_rshift_data;
  reg __mul_13_stream_ivalid_1;
  reg __mul_13_stream_ivalid_2;
  reg __mul_13_stream_ivalid_3;
  reg __mul_13_stream_ivalid_4;
  reg __mul_13_stream_ivalid_5;
  reg __mul_13_stream_ivalid_6;
  reg __mul_13_stream_ivalid_7;
  reg __mul_13_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_244;
  reg [5-1:0] _minus_data_246;
  reg [1-1:0] _greatereq_data_257;
  reg signed [16-1:0] __delay_data_816__variable_241;
  reg signed [16-1:0] __delay_data_819__variable_242;
  reg [5-1:0] __delay_data_822__variable_243;
  reg signed [34-1:0] _sll_data_248;
  reg [1-1:0] __delay_data_813_greaterthan_244;
  reg [1-1:0] __delay_data_814_greatereq_257;
  reg signed [16-1:0] __delay_data_817__delay_816__variable_241;
  reg signed [16-1:0] __delay_data_820__delay_819__variable_242;
  reg [5-1:0] __delay_data_823__delay_822__variable_243;
  reg signed [32-1:0] _cond_data_254;
  reg [1-1:0] __delay_data_815__delay_814_greatereq_257;
  reg signed [16-1:0] __delay_data_818__delay_817__delay_816__variable_241;
  reg signed [16-1:0] __delay_data_821__delay_820__delay_819__variable_242;
  reg [5-1:0] __delay_data_824__delay_823__delay_822__variable_243;
  wire signed [16-1:0] _uminus_data_256;
  assign _uminus_data_256 = -_cond_data_254;
  wire signed [16-1:0] _cond_data_259;
  assign _cond_data_259 = (__delay_data_815__delay_814_greatereq_257)? _cond_data_254 : _uminus_data_256;
  wire signed [32-1:0] __muladd_madd_odata_260;
  reg signed [32-1:0] __muladd_madd_odata_reg_260;
  wire signed [32-1:0] __muladd_data_260;
  assign __muladd_data_260 = __muladd_madd_odata_reg_260;
  wire __muladd_madd_update_260;
  assign __muladd_madd_update_260 = _mul_13_stream_oready;

  madd_5
  __muladd_madd_260
  (
    .CLK(CLK),
    .update(__muladd_madd_update_260),
    .a(__delay_data_818__delay_817__delay_816__variable_241),
    .b(__delay_data_821__delay_820__delay_819__variable_242),
    .c(_cond_data_259),
    .d(__muladd_madd_odata_260)
  );

  reg [5-1:0] __delay_data_825__delay_824__delay_823____variable_243;
  reg [5-1:0] __delay_data_826__delay_825__delay_824____variable_243;
  reg [5-1:0] __delay_data_827__delay_826__delay_825____variable_243;
  reg [5-1:0] __delay_data_828__delay_827__delay_826____variable_243;
  reg signed [32-1:0] _sra_data_261;
  wire signed [32-1:0] mul_13_z_data;
  assign mul_13_z_data = _sra_data_261;
  wire signed [16-1:0] mul_14_x_data;
  wire signed [16-1:0] mul_14_y_data;
  wire [5-1:0] mul_14_rshift_data;
  reg __mul_14_stream_ivalid_1;
  reg __mul_14_stream_ivalid_2;
  reg __mul_14_stream_ivalid_3;
  reg __mul_14_stream_ivalid_4;
  reg __mul_14_stream_ivalid_5;
  reg __mul_14_stream_ivalid_6;
  reg __mul_14_stream_ivalid_7;
  reg __mul_14_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_265;
  reg [5-1:0] _minus_data_267;
  reg [1-1:0] _greatereq_data_278;
  reg signed [16-1:0] __delay_data_835__variable_262;
  reg signed [16-1:0] __delay_data_838__variable_263;
  reg [5-1:0] __delay_data_841__variable_264;
  reg signed [34-1:0] _sll_data_269;
  reg [1-1:0] __delay_data_832_greaterthan_265;
  reg [1-1:0] __delay_data_833_greatereq_278;
  reg signed [16-1:0] __delay_data_836__delay_835__variable_262;
  reg signed [16-1:0] __delay_data_839__delay_838__variable_263;
  reg [5-1:0] __delay_data_842__delay_841__variable_264;
  reg signed [32-1:0] _cond_data_275;
  reg [1-1:0] __delay_data_834__delay_833_greatereq_278;
  reg signed [16-1:0] __delay_data_837__delay_836__delay_835__variable_262;
  reg signed [16-1:0] __delay_data_840__delay_839__delay_838__variable_263;
  reg [5-1:0] __delay_data_843__delay_842__delay_841__variable_264;
  wire signed [16-1:0] _uminus_data_277;
  assign _uminus_data_277 = -_cond_data_275;
  wire signed [16-1:0] _cond_data_280;
  assign _cond_data_280 = (__delay_data_834__delay_833_greatereq_278)? _cond_data_275 : _uminus_data_277;
  wire signed [32-1:0] __muladd_madd_odata_281;
  reg signed [32-1:0] __muladd_madd_odata_reg_281;
  wire signed [32-1:0] __muladd_data_281;
  assign __muladd_data_281 = __muladd_madd_odata_reg_281;
  wire __muladd_madd_update_281;
  assign __muladd_madd_update_281 = _mul_14_stream_oready;

  madd_6
  __muladd_madd_281
  (
    .CLK(CLK),
    .update(__muladd_madd_update_281),
    .a(__delay_data_837__delay_836__delay_835__variable_262),
    .b(__delay_data_840__delay_839__delay_838__variable_263),
    .c(_cond_data_280),
    .d(__muladd_madd_odata_281)
  );

  reg [5-1:0] __delay_data_844__delay_843__delay_842____variable_264;
  reg [5-1:0] __delay_data_845__delay_844__delay_843____variable_264;
  reg [5-1:0] __delay_data_846__delay_845__delay_844____variable_264;
  reg [5-1:0] __delay_data_847__delay_846__delay_845____variable_264;
  reg signed [32-1:0] _sra_data_282;
  wire signed [32-1:0] mul_14_z_data;
  assign mul_14_z_data = _sra_data_282;
  wire signed [16-1:0] mul_15_x_data;
  wire signed [16-1:0] mul_15_y_data;
  wire [5-1:0] mul_15_rshift_data;
  reg __mul_15_stream_ivalid_1;
  reg __mul_15_stream_ivalid_2;
  reg __mul_15_stream_ivalid_3;
  reg __mul_15_stream_ivalid_4;
  reg __mul_15_stream_ivalid_5;
  reg __mul_15_stream_ivalid_6;
  reg __mul_15_stream_ivalid_7;
  reg __mul_15_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_286;
  reg [5-1:0] _minus_data_288;
  reg [1-1:0] _greatereq_data_299;
  reg signed [16-1:0] __delay_data_854__variable_283;
  reg signed [16-1:0] __delay_data_857__variable_284;
  reg [5-1:0] __delay_data_860__variable_285;
  reg signed [34-1:0] _sll_data_290;
  reg [1-1:0] __delay_data_851_greaterthan_286;
  reg [1-1:0] __delay_data_852_greatereq_299;
  reg signed [16-1:0] __delay_data_855__delay_854__variable_283;
  reg signed [16-1:0] __delay_data_858__delay_857__variable_284;
  reg [5-1:0] __delay_data_861__delay_860__variable_285;
  reg signed [32-1:0] _cond_data_296;
  reg [1-1:0] __delay_data_853__delay_852_greatereq_299;
  reg signed [16-1:0] __delay_data_856__delay_855__delay_854__variable_283;
  reg signed [16-1:0] __delay_data_859__delay_858__delay_857__variable_284;
  reg [5-1:0] __delay_data_862__delay_861__delay_860__variable_285;
  wire signed [16-1:0] _uminus_data_298;
  assign _uminus_data_298 = -_cond_data_296;
  wire signed [16-1:0] _cond_data_301;
  assign _cond_data_301 = (__delay_data_853__delay_852_greatereq_299)? _cond_data_296 : _uminus_data_298;
  wire signed [32-1:0] __muladd_madd_odata_302;
  reg signed [32-1:0] __muladd_madd_odata_reg_302;
  wire signed [32-1:0] __muladd_data_302;
  assign __muladd_data_302 = __muladd_madd_odata_reg_302;
  wire __muladd_madd_update_302;
  assign __muladd_madd_update_302 = _mul_15_stream_oready;

  madd_7
  __muladd_madd_302
  (
    .CLK(CLK),
    .update(__muladd_madd_update_302),
    .a(__delay_data_856__delay_855__delay_854__variable_283),
    .b(__delay_data_859__delay_858__delay_857__variable_284),
    .c(_cond_data_301),
    .d(__muladd_madd_odata_302)
  );

  reg [5-1:0] __delay_data_863__delay_862__delay_861____variable_285;
  reg [5-1:0] __delay_data_864__delay_863__delay_862____variable_285;
  reg [5-1:0] __delay_data_865__delay_864__delay_863____variable_285;
  reg [5-1:0] __delay_data_866__delay_865__delay_864____variable_285;
  reg signed [32-1:0] _sra_data_303;
  wire signed [32-1:0] mul_15_z_data;
  assign mul_15_z_data = _sra_data_303;
  wire signed [16-1:0] mul_16_x_data;
  wire signed [16-1:0] mul_16_y_data;
  wire [5-1:0] mul_16_rshift_data;
  reg __mul_16_stream_ivalid_1;
  reg __mul_16_stream_ivalid_2;
  reg __mul_16_stream_ivalid_3;
  reg __mul_16_stream_ivalid_4;
  reg __mul_16_stream_ivalid_5;
  reg __mul_16_stream_ivalid_6;
  reg __mul_16_stream_ivalid_7;
  reg __mul_16_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_307;
  reg [5-1:0] _minus_data_309;
  reg [1-1:0] _greatereq_data_320;
  reg signed [16-1:0] __delay_data_873__variable_304;
  reg signed [16-1:0] __delay_data_876__variable_305;
  reg [5-1:0] __delay_data_879__variable_306;
  reg signed [34-1:0] _sll_data_311;
  reg [1-1:0] __delay_data_870_greaterthan_307;
  reg [1-1:0] __delay_data_871_greatereq_320;
  reg signed [16-1:0] __delay_data_874__delay_873__variable_304;
  reg signed [16-1:0] __delay_data_877__delay_876__variable_305;
  reg [5-1:0] __delay_data_880__delay_879__variable_306;
  reg signed [32-1:0] _cond_data_317;
  reg [1-1:0] __delay_data_872__delay_871_greatereq_320;
  reg signed [16-1:0] __delay_data_875__delay_874__delay_873__variable_304;
  reg signed [16-1:0] __delay_data_878__delay_877__delay_876__variable_305;
  reg [5-1:0] __delay_data_881__delay_880__delay_879__variable_306;
  wire signed [16-1:0] _uminus_data_319;
  assign _uminus_data_319 = -_cond_data_317;
  wire signed [16-1:0] _cond_data_322;
  assign _cond_data_322 = (__delay_data_872__delay_871_greatereq_320)? _cond_data_317 : _uminus_data_319;
  wire signed [32-1:0] __muladd_madd_odata_323;
  reg signed [32-1:0] __muladd_madd_odata_reg_323;
  wire signed [32-1:0] __muladd_data_323;
  assign __muladd_data_323 = __muladd_madd_odata_reg_323;
  wire __muladd_madd_update_323;
  assign __muladd_madd_update_323 = _mul_16_stream_oready;

  madd_8
  __muladd_madd_323
  (
    .CLK(CLK),
    .update(__muladd_madd_update_323),
    .a(__delay_data_875__delay_874__delay_873__variable_304),
    .b(__delay_data_878__delay_877__delay_876__variable_305),
    .c(_cond_data_322),
    .d(__muladd_madd_odata_323)
  );

  reg [5-1:0] __delay_data_882__delay_881__delay_880____variable_306;
  reg [5-1:0] __delay_data_883__delay_882__delay_881____variable_306;
  reg [5-1:0] __delay_data_884__delay_883__delay_882____variable_306;
  reg [5-1:0] __delay_data_885__delay_884__delay_883____variable_306;
  reg signed [32-1:0] _sra_data_324;
  wire signed [32-1:0] mul_16_z_data;
  assign mul_16_z_data = _sra_data_324;
  wire signed [64-1:0] add_tree_5_var0_data;
  wire signed [64-1:0] add_tree_5_var1_data;
  wire signed [64-1:0] add_tree_5_var2_data;
  wire signed [64-1:0] add_tree_5_var3_data;
  wire signed [64-1:0] add_tree_5_var4_data;
  wire signed [64-1:0] add_tree_5_var5_data;
  wire signed [64-1:0] add_tree_5_var6_data;
  wire signed [64-1:0] add_tree_5_var7_data;
  wire signed [64-1:0] add_tree_5_var8_data;
  reg __add_tree_5_stream_ivalid_1;
  reg __add_tree_5_stream_ivalid_2;
  reg signed [64-1:0] __plusn_data_64;
  reg signed [64-1:0] __plusn_data_65;
  reg signed [64-1:0] __plusn_data_66;
  reg signed [64-1:0] __plusn_data_67;
  wire signed [64-1:0] add_tree_5_sum_data;
  assign add_tree_5_sum_data = __plusn_data_67;
  wire signed [64-1:0] acc_0_x_data;
  wire [7-1:0] acc_0_rshift_data;
  wire [32-1:0] acc_0_size_data;
  wire [1-1:0] acc_0__reduce_reset_data;
  reg __acc_0_stream_ivalid_1;
  reg __acc_0_stream_ivalid_2;
  reg __acc_0_stream_ivalid_3;
  reg __acc_0_stream_ivalid_4;
  reg __acc_0_stream_ivalid_5;
  reg [1-1:0] _greaterthan_data_3;
  reg [7-1:0] _minus_data_5;
  reg signed [64-1:0] _reduceadd_data_16;
  reg [33-1:0] _reduceadd_count_16;
  reg _reduceadd_prev_count_max_16;
  wire _reduceadd_reset_cond_16;
  assign _reduceadd_reset_cond_16 = acc_0__reduce_reset_data || _reduceadd_prev_count_max_16;
  wire [33-1:0] _reduceadd_current_count_16;
  assign _reduceadd_current_count_16 = (_reduceadd_reset_cond_16)? 0 : _reduceadd_count_16;
  wire signed [64-1:0] _reduceadd_current_data_16;
  assign _reduceadd_current_data_16 = (_reduceadd_reset_cond_16)? 1'sd0 : _reduceadd_data_16;
  reg [1-1:0] _pulse_data_18;
  reg [33-1:0] _pulse_count_18;
  reg _pulse_prev_count_max_18;
  wire _pulse_reset_cond_18;
  assign _pulse_reset_cond_18 = acc_0__reduce_reset_data || _pulse_prev_count_max_18;
  wire [33-1:0] _pulse_current_count_18;
  assign _pulse_current_count_18 = (_pulse_reset_cond_18)? 0 : _pulse_count_18;
  wire [1-1:0] _pulse_current_data_18;
  assign _pulse_current_data_18 = (_pulse_reset_cond_18)? 1'sd0 : _pulse_data_18;
  reg [7-1:0] __delay_data_894__variable_1;
  reg signed [130-1:0] _sll_data_7;
  reg [1-1:0] __delay_data_891_greaterthan_3;
  reg signed [64-1:0] __delay_data_892_reduceadd_16;
  reg [7-1:0] __delay_data_895__delay_894__variable_1;
  reg [1-1:0] __delay_data_898_pulse_18;
  reg signed [64-1:0] _cond_data_13;
  reg signed [64-1:0] __delay_data_893__delay_892_reduceadd_16;
  reg [7-1:0] __delay_data_896__delay_895__delay_894__variable_1;
  reg [1-1:0] __delay_data_899__delay_898_pulse_18;
  reg signed [64-1:0] _plus_data_20;
  reg [7-1:0] __delay_data_897__delay_896__delay_895__delay_894__variable_1;
  reg [1-1:0] __delay_data_900__delay_899__delay_898_pulse_18;
  reg signed [64-1:0] _sra_data_21;
  reg [1-1:0] __delay_data_901__delay_900__delay_899__delay_898_pulse_18;
  wire signed [64-1:0] acc_0_sum_data;
  assign acc_0_sum_data = _sra_data_21;
  wire [1-1:0] acc_0_valid_data;
  assign acc_0_valid_data = __delay_data_901__delay_900__delay_899__delay_898_pulse_18;
  wire signed [64-1:0] mul_rshift_round_clip_6_x_data;
  wire signed [16-1:0] mul_rshift_round_clip_6_y_data;
  wire [7-1:0] mul_rshift_round_clip_6_rshift_data;
  reg __mul_rshift_round_clip_6_stream_ivalid_1;
  reg __mul_rshift_round_clip_6_stream_ivalid_2;
  reg __mul_rshift_round_clip_6_stream_ivalid_3;
  reg __mul_rshift_round_clip_6_stream_ivalid_4;
  reg __mul_rshift_round_clip_6_stream_ivalid_5;
  reg __mul_rshift_round_clip_6_stream_ivalid_6;
  reg __mul_rshift_round_clip_6_stream_ivalid_7;
  reg __mul_rshift_round_clip_6_stream_ivalid_8;
  wire signed [80-1:0] _times_mul_odata_71;
  reg signed [80-1:0] _times_mul_odata_reg_71;
  wire signed [80-1:0] _times_data_71;
  assign _times_data_71 = _times_mul_odata_reg_71;
  wire _times_mul_update_71;
  assign _times_mul_update_71 = _mul_rshift_round_clip_6_stream_oready;

  multiplier_0
  _times_mul_71
  (
    .CLK(CLK),
    .update(_times_mul_update_71),
    .a(mul_rshift_round_clip_6_x_data),
    .b(mul_rshift_round_clip_6_y_data),
    .c(_times_mul_odata_71)
  );

  wire [7-1:0] _minus_data_74;
  assign _minus_data_74 = mul_rshift_round_clip_6_rshift_data - 2'sd1;
  wire signed [130-1:0] _sll_data_77;
  assign _sll_data_77 = 2'sd1 << _minus_data_74;
  wire [1-1:0] _eq_data_89;
  assign _eq_data_89 = mul_rshift_round_clip_6_rshift_data == 1'sd0;
  reg signed [130-1:0] __delay_data_907_sll_77;
  reg [7-1:0] __delay_data_911__variable_70;
  reg [1-1:0] __delay_data_915_eq_89;
  reg signed [130-1:0] __delay_data_908__delay_907_sll_77;
  reg [7-1:0] __delay_data_912__delay_911__variable_70;
  reg [1-1:0] __delay_data_916__delay_915_eq_89;
  reg signed [130-1:0] __delay_data_909__delay_908__delay_907_sll_77;
  reg [7-1:0] __delay_data_913__delay_912__delay_911__variable_70;
  reg [1-1:0] __delay_data_917__delay_916__delay_915_eq_89;
  reg signed [130-1:0] __delay_data_910__delay_909__delay_908__delay_907_sll_77;
  reg [7-1:0] __delay_data_914__delay_913__delay_912__delay_911__variable_70;
  reg [1-1:0] __delay_data_918__delay_917__delay_916__delay_915_eq_89;
  wire [1-1:0] _pointer_data_72;
  assign _pointer_data_72 = _times_data_71[8'sd79];
  wire signed [2-1:0] _cond_data_84;
  assign _cond_data_84 = (_pointer_data_72)? -2'sd1 : 1'sd0;
  wire signed [81-1:0] _plus_data_85;
  assign _plus_data_85 = _times_data_71 + __delay_data_910__delay_909__delay_908__delay_907_sll_77;
  wire signed [81-1:0] _plus_data_86;
  assign _plus_data_86 = _plus_data_85 + _cond_data_84;
  wire signed [80-1:0] _sra_data_87;
  assign _sra_data_87 = _plus_data_86 >>> __delay_data_914__delay_913__delay_912__delay_911__variable_70;
  reg signed [80-1:0] _cond_data_90;
  reg [1-1:0] _greaterthan_data_91;
  reg [1-1:0] _lessthan_data_95;
  reg [1-1:0] _greatereq_data_99;
  reg signed [80-1:0] __delay_data_919_cond_90;
  reg signed [80-1:0] _cond_data_93;
  reg signed [80-1:0] _cond_data_97;
  reg [1-1:0] __delay_data_920_greatereq_99;
  reg signed [16-1:0] _cond_data_101;
  wire signed [16-1:0] mul_rshift_round_clip_6_z_data;
  assign mul_rshift_round_clip_6_z_data = _cond_data_101;
  reg [33-1:0] _stream_conv2d_4_sink_50_sink_count;
  reg [5-1:0] _stream_conv2d_4_sink_50_sink_mode;
  reg [16-1:0] _stream_conv2d_4_sink_50_sink_generator_id;
  reg [32-1:0] _stream_conv2d_4_sink_50_sink_offset;
  reg [33-1:0] _stream_conv2d_4_sink_50_sink_size;
  reg [32-1:0] _stream_conv2d_4_sink_50_sink_stride;
  reg [32-1:0] _stream_conv2d_4_sink_50_sink_offset_buf;
  reg [33-1:0] _stream_conv2d_4_sink_50_sink_size_buf;
  reg [32-1:0] _stream_conv2d_4_sink_50_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_4_sink_50_sink_sel;
  reg [32-1:0] _stream_conv2d_4_sink_50_sink_waddr;
  reg _stream_conv2d_4_sink_50_sink_wenable;
  reg [16-1:0] _stream_conv2d_4_sink_50_sink_wdata;
  reg _stream_conv2d_4_sink_50_sink_fifo_enq;
  reg [16-1:0] _stream_conv2d_4_sink_50_sink_fifo_wdata;
  reg [16-1:0] _stream_conv2d_4_sink_50_sink_immediate;
  reg [33-1:0] _stream_conv2d_4_sink_51_sink_count;
  reg [5-1:0] _stream_conv2d_4_sink_51_sink_mode;
  reg [16-1:0] _stream_conv2d_4_sink_51_sink_generator_id;
  reg [32-1:0] _stream_conv2d_4_sink_51_sink_offset;
  reg [33-1:0] _stream_conv2d_4_sink_51_sink_size;
  reg [32-1:0] _stream_conv2d_4_sink_51_sink_stride;
  reg [32-1:0] _stream_conv2d_4_sink_51_sink_offset_buf;
  reg [33-1:0] _stream_conv2d_4_sink_51_sink_size_buf;
  reg [32-1:0] _stream_conv2d_4_sink_51_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_4_sink_51_sink_sel;
  reg [32-1:0] _stream_conv2d_4_sink_51_sink_waddr;
  reg _stream_conv2d_4_sink_51_sink_wenable;
  reg [1-1:0] _stream_conv2d_4_sink_51_sink_wdata;
  reg _stream_conv2d_4_sink_51_sink_fifo_enq;
  reg [1-1:0] _stream_conv2d_4_sink_51_sink_fifo_wdata;
  reg [1-1:0] _stream_conv2d_4_sink_51_sink_immediate;
  reg _stream_max_pool_serial_6_stream_ivalid;
  wire _stream_max_pool_serial_6_stream_oready;
  wire _stream_max_pool_serial_6_stream_internal_oready;
  assign _stream_max_pool_serial_6_stream_oready = _stream_max_pool_serial_6_stream_internal_oready;
  reg [32-1:0] _stream_max_pool_serial_6_fsm;
  localparam _stream_max_pool_serial_6_fsm_init = 0;
  wire _stream_max_pool_serial_6_run_flag;
  reg _stream_max_pool_serial_6_source_start;
  wire _stream_max_pool_serial_6_source_stop;
  reg _stream_max_pool_serial_6_source_busy;
  wire _stream_max_pool_serial_6_sink_start;
  wire _stream_max_pool_serial_6_sink_stop;
  wire _stream_max_pool_serial_6_sink_busy;
  wire _stream_max_pool_serial_6_busy;
  reg _stream_max_pool_serial_6_busy_reg;
  wire _stream_max_pool_serial_6_is_root;
  assign _stream_max_pool_serial_6_is_root = 1;
  reg [3-1:0] _stream_max_pool_serial_6_parameter_0_next_parameter_data;
  reg _stream_max_pool_serial_6_source_1_idle;
  reg [33-1:0] _stream_max_pool_serial_6_source_1_source_count;
  reg [5-1:0] _stream_max_pool_serial_6_source_1_source_mode;
  reg [16-1:0] _stream_max_pool_serial_6_source_1_source_generator_id;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_offset;
  reg [33-1:0] _stream_max_pool_serial_6_source_1_source_size;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_stride;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_6_source_1_source_size_buf;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_6_source_1_source_sel;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_ram_raddr;
  reg _stream_max_pool_serial_6_source_1_source_ram_renable;
  wire [32-1:0] _stream_max_pool_serial_6_source_1_source_ram_rdata;
  reg _stream_max_pool_serial_6_source_1_source_fifo_deq;
  wire [32-1:0] _stream_max_pool_serial_6_source_1_source_fifo_rdata;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_empty_data;
  reg [4-1:0] _stream_max_pool_serial_6_parameter_2_next_parameter_data;
  wire signed [16-1:0] _reduce_max_17_x_data;
  wire [32-1:0] _reduce_max_17_size_data;
  wire [1-1:0] _reduce_max_17__reduce_reset_data;
  reg ___reduce_max_17_stream_ivalid_1;
  reg signed [16-1:0] _reducemax_data_328;
  reg [33-1:0] _reducemax_count_328;
  reg _reducemax_prev_count_max_328;
  wire _reducemax_reset_cond_328;
  assign _reducemax_reset_cond_328 = _reduce_max_17__reduce_reset_data || _reducemax_prev_count_max_328;
  wire [33-1:0] _reducemax_current_count_328;
  assign _reducemax_current_count_328 = (_reducemax_reset_cond_328)? 0 : _reducemax_count_328;
  wire signed [16-1:0] _reducemax_current_data_328;
  assign _reducemax_current_data_328 = (_reducemax_reset_cond_328)? -17'sd32768 : _reducemax_data_328;
  reg [1-1:0] _pulse_data_330;
  reg [33-1:0] _pulse_count_330;
  reg _pulse_prev_count_max_330;
  wire _pulse_reset_cond_330;
  assign _pulse_reset_cond_330 = _reduce_max_17__reduce_reset_data || _pulse_prev_count_max_330;
  wire [33-1:0] _pulse_current_count_330;
  assign _pulse_current_count_330 = (_pulse_reset_cond_330)? 0 : _pulse_count_330;
  wire [1-1:0] _pulse_current_data_330;
  assign _pulse_current_data_330 = (_pulse_reset_cond_330)? 1'sd0 : _pulse_data_330;
  wire signed [16-1:0] _reduce_max_17_data_data;
  assign _reduce_max_17_data_data = _reducemax_data_328;
  wire [1-1:0] _reduce_max_17_valid_data;
  assign _reduce_max_17_valid_data = _pulse_data_330;
  wire signed [16-1:0] _reduce_max_18_x_data;
  wire [32-1:0] _reduce_max_18_size_data;
  wire [1-1:0] _reduce_max_18__reduce_reset_data;
  reg ___reduce_max_18_stream_ivalid_1;
  reg signed [16-1:0] _reducemax_data_335;
  reg [33-1:0] _reducemax_count_335;
  reg _reducemax_prev_count_max_335;
  wire _reducemax_reset_cond_335;
  assign _reducemax_reset_cond_335 = _reduce_max_18__reduce_reset_data || _reducemax_prev_count_max_335;
  wire [33-1:0] _reducemax_current_count_335;
  assign _reducemax_current_count_335 = (_reducemax_reset_cond_335)? 0 : _reducemax_count_335;
  wire signed [16-1:0] _reducemax_current_data_335;
  assign _reducemax_current_data_335 = (_reducemax_reset_cond_335)? -17'sd32768 : _reducemax_data_335;
  reg [1-1:0] _pulse_data_337;
  reg [33-1:0] _pulse_count_337;
  reg _pulse_prev_count_max_337;
  wire _pulse_reset_cond_337;
  assign _pulse_reset_cond_337 = _reduce_max_18__reduce_reset_data || _pulse_prev_count_max_337;
  wire [33-1:0] _pulse_current_count_337;
  assign _pulse_current_count_337 = (_pulse_reset_cond_337)? 0 : _pulse_count_337;
  wire [1-1:0] _pulse_current_data_337;
  assign _pulse_current_data_337 = (_pulse_reset_cond_337)? 1'sd0 : _pulse_data_337;
  wire signed [16-1:0] _reduce_max_18_data_data;
  assign _reduce_max_18_data_data = _reducemax_data_335;
  wire [1-1:0] _reduce_max_18_valid_data;
  assign _reduce_max_18_valid_data = _pulse_data_337;
  reg [33-1:0] _stream_max_pool_serial_6_sink_6_sink_count;
  reg [5-1:0] _stream_max_pool_serial_6_sink_6_sink_mode;
  reg [16-1:0] _stream_max_pool_serial_6_sink_6_sink_generator_id;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_offset;
  reg [33-1:0] _stream_max_pool_serial_6_sink_6_sink_size;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_stride;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_6_sink_6_sink_size_buf;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_6_sink_6_sink_sel;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_waddr;
  reg _stream_max_pool_serial_6_sink_6_sink_wenable;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_wdata;
  reg _stream_max_pool_serial_6_sink_6_sink_fifo_enq;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_fifo_wdata;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_immediate;
  reg [33-1:0] _stream_max_pool_serial_6_sink_7_sink_count;
  reg [5-1:0] _stream_max_pool_serial_6_sink_7_sink_mode;
  reg [16-1:0] _stream_max_pool_serial_6_sink_7_sink_generator_id;
  reg [32-1:0] _stream_max_pool_serial_6_sink_7_sink_offset;
  reg [33-1:0] _stream_max_pool_serial_6_sink_7_sink_size;
  reg [32-1:0] _stream_max_pool_serial_6_sink_7_sink_stride;
  reg [32-1:0] _stream_max_pool_serial_6_sink_7_sink_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_6_sink_7_sink_size_buf;
  reg [32-1:0] _stream_max_pool_serial_6_sink_7_sink_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_6_sink_7_sink_sel;
  reg [32-1:0] _stream_max_pool_serial_6_sink_7_sink_waddr;
  reg _stream_max_pool_serial_6_sink_7_sink_wenable;
  reg [1-1:0] _stream_max_pool_serial_6_sink_7_sink_wdata;
  reg _stream_max_pool_serial_6_sink_7_sink_fifo_enq;
  reg [1-1:0] _stream_max_pool_serial_6_sink_7_sink_fifo_wdata;
  reg [1-1:0] _stream_max_pool_serial_6_sink_7_sink_immediate;
  reg _stream_matmul_23_stream_ivalid;
  wire _stream_matmul_23_stream_oready;
  wire _stream_matmul_23_stream_internal_oready;
  assign _stream_matmul_23_stream_oready = _stream_matmul_23_stream_internal_oready;
  reg [32-1:0] _stream_matmul_23_fsm;
  localparam _stream_matmul_23_fsm_init = 0;
  wire _stream_matmul_23_run_flag;
  reg _stream_matmul_23_source_start;
  wire _stream_matmul_23_source_stop;
  reg _stream_matmul_23_source_busy;
  wire _stream_matmul_23_sink_start;
  wire _stream_matmul_23_sink_stop;
  wire _stream_matmul_23_sink_busy;
  wire _stream_matmul_23_busy;
  reg _stream_matmul_23_busy_reg;
  wire _stream_matmul_23_is_root;
  assign _stream_matmul_23_is_root = 1;
  reg [13-1:0] _stream_matmul_23_parameter_0_next_parameter_data;
  reg [1-1:0] _stream_matmul_23_parameter_1_next_parameter_data;
  reg [1-1:0] _stream_matmul_23_parameter_2_next_parameter_data;
  reg [1-1:0] _stream_matmul_23_parameter_3_next_parameter_data;
  reg [1-1:0] _stream_matmul_23_parameter_4_next_parameter_data;
  reg [1-1:0] _stream_matmul_23_parameter_6_next_parameter_data;
  reg _stream_matmul_23_source_7_idle;
  reg [33-1:0] _stream_matmul_23_source_7_source_count;
  reg [5-1:0] _stream_matmul_23_source_7_source_mode;
  reg [16-1:0] _stream_matmul_23_source_7_source_generator_id;
  reg [32-1:0] _stream_matmul_23_source_7_source_offset;
  reg [33-1:0] _stream_matmul_23_source_7_source_size;
  reg [32-1:0] _stream_matmul_23_source_7_source_stride;
  reg [32-1:0] _stream_matmul_23_source_7_source_offset_buf;
  reg [33-1:0] _stream_matmul_23_source_7_source_size_buf;
  reg [32-1:0] _stream_matmul_23_source_7_source_stride_buf;
  reg [8-1:0] _stream_matmul_23_source_7_source_sel;
  reg [32-1:0] _stream_matmul_23_source_7_source_ram_raddr;
  reg _stream_matmul_23_source_7_source_ram_renable;
  wire [16-1:0] _stream_matmul_23_source_7_source_ram_rdata;
  reg _stream_matmul_23_source_7_source_fifo_deq;
  wire [16-1:0] _stream_matmul_23_source_7_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_23_source_7_source_empty_data;
  reg [1-1:0] _stream_matmul_23_parameter_8_next_parameter_data;
  reg _stream_matmul_23_source_9_idle;
  reg [33-1:0] _stream_matmul_23_source_9_source_count;
  reg [5-1:0] _stream_matmul_23_source_9_source_mode;
  reg [16-1:0] _stream_matmul_23_source_9_source_generator_id;
  reg [32-1:0] _stream_matmul_23_source_9_source_offset;
  reg [33-1:0] _stream_matmul_23_source_9_source_size;
  reg [32-1:0] _stream_matmul_23_source_9_source_stride;
  reg [32-1:0] _stream_matmul_23_source_9_source_offset_buf;
  reg [33-1:0] _stream_matmul_23_source_9_source_size_buf;
  reg [32-1:0] _stream_matmul_23_source_9_source_stride_buf;
  reg [8-1:0] _stream_matmul_23_source_9_source_sel;
  reg [32-1:0] _stream_matmul_23_source_9_source_ram_raddr;
  reg _stream_matmul_23_source_9_source_ram_renable;
  wire [16-1:0] _stream_matmul_23_source_9_source_ram_rdata;
  reg _stream_matmul_23_source_9_source_fifo_deq;
  wire [16-1:0] _stream_matmul_23_source_9_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_23_source_9_source_empty_data;
  reg [1-1:0] _stream_matmul_23_parameter_10_next_parameter_data;
  reg _stream_matmul_23_source_11_idle;
  reg [33-1:0] _stream_matmul_23_source_11_source_count;
  reg [5-1:0] _stream_matmul_23_source_11_source_mode;
  reg [16-1:0] _stream_matmul_23_source_11_source_generator_id;
  reg [32-1:0] _stream_matmul_23_source_11_source_offset;
  reg [33-1:0] _stream_matmul_23_source_11_source_size;
  reg [32-1:0] _stream_matmul_23_source_11_source_stride;
  reg [32-1:0] _stream_matmul_23_source_11_source_offset_buf;
  reg [33-1:0] _stream_matmul_23_source_11_source_size_buf;
  reg [32-1:0] _stream_matmul_23_source_11_source_stride_buf;
  reg [8-1:0] _stream_matmul_23_source_11_source_sel;
  reg [32-1:0] _stream_matmul_23_source_11_source_ram_raddr;
  reg _stream_matmul_23_source_11_source_ram_renable;
  wire [16-1:0] _stream_matmul_23_source_11_source_ram_rdata;
  reg _stream_matmul_23_source_11_source_fifo_deq;
  wire [16-1:0] _stream_matmul_23_source_11_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_23_source_11_source_empty_data;
  reg [1-1:0] _stream_matmul_23_parameter_12_next_parameter_data;
  reg _stream_matmul_23_source_13_idle;
  reg [33-1:0] _stream_matmul_23_source_13_source_count;
  reg [5-1:0] _stream_matmul_23_source_13_source_mode;
  reg [16-1:0] _stream_matmul_23_source_13_source_generator_id;
  reg [32-1:0] _stream_matmul_23_source_13_source_offset;
  reg [33-1:0] _stream_matmul_23_source_13_source_size;
  reg [32-1:0] _stream_matmul_23_source_13_source_stride;
  reg [32-1:0] _stream_matmul_23_source_13_source_offset_buf;
  reg [33-1:0] _stream_matmul_23_source_13_source_size_buf;
  reg [32-1:0] _stream_matmul_23_source_13_source_stride_buf;
  reg [8-1:0] _stream_matmul_23_source_13_source_sel;
  reg [32-1:0] _stream_matmul_23_source_13_source_ram_raddr;
  reg _stream_matmul_23_source_13_source_ram_renable;
  wire [16-1:0] _stream_matmul_23_source_13_source_ram_rdata;
  reg _stream_matmul_23_source_13_source_fifo_deq;
  wire [16-1:0] _stream_matmul_23_source_13_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_23_source_13_source_empty_data;
  reg [1-1:0] _stream_matmul_23_parameter_14_next_parameter_data;
  reg _stream_matmul_23_source_15_idle;
  reg [33-1:0] _stream_matmul_23_source_15_source_count;
  reg [5-1:0] _stream_matmul_23_source_15_source_mode;
  reg [16-1:0] _stream_matmul_23_source_15_source_generator_id;
  reg [32-1:0] _stream_matmul_23_source_15_source_offset;
  reg [33-1:0] _stream_matmul_23_source_15_source_size;
  reg [32-1:0] _stream_matmul_23_source_15_source_stride;
  reg [32-1:0] _stream_matmul_23_source_15_source_offset_buf;
  reg [33-1:0] _stream_matmul_23_source_15_source_size_buf;
  reg [32-1:0] _stream_matmul_23_source_15_source_stride_buf;
  reg [8-1:0] _stream_matmul_23_source_15_source_sel;
  reg [32-1:0] _stream_matmul_23_source_15_source_ram_raddr;
  reg _stream_matmul_23_source_15_source_ram_renable;
  wire [16-1:0] _stream_matmul_23_source_15_source_ram_rdata;
  reg _stream_matmul_23_source_15_source_fifo_deq;
  wire [16-1:0] _stream_matmul_23_source_15_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_23_source_15_source_empty_data;
  reg [1-1:0] _stream_matmul_23_parameter_16_next_parameter_data;
  reg [1-1:0] _stream_matmul_23_parameter_17_next_parameter_data;
  reg [1-1:0] _stream_matmul_23_parameter_18_next_parameter_data;
  reg [1-1:0] _stream_matmul_23_parameter_19_next_parameter_data;
  reg _stream_matmul_23_source_20_idle;
  reg [33-1:0] _stream_matmul_23_source_20_source_count;
  reg [5-1:0] _stream_matmul_23_source_20_source_mode;
  reg [16-1:0] _stream_matmul_23_source_20_source_generator_id;
  reg [32-1:0] _stream_matmul_23_source_20_source_offset;
  reg [33-1:0] _stream_matmul_23_source_20_source_size;
  reg [32-1:0] _stream_matmul_23_source_20_source_stride;
  reg [32-1:0] _stream_matmul_23_source_20_source_offset_buf;
  reg [33-1:0] _stream_matmul_23_source_20_source_size_buf;
  reg [32-1:0] _stream_matmul_23_source_20_source_stride_buf;
  reg [8-1:0] _stream_matmul_23_source_20_source_sel;
  reg [32-1:0] _stream_matmul_23_source_20_source_ram_raddr;
  reg _stream_matmul_23_source_20_source_ram_renable;
  wire [16-1:0] _stream_matmul_23_source_20_source_ram_rdata;
  reg _stream_matmul_23_source_20_source_fifo_deq;
  wire [16-1:0] _stream_matmul_23_source_20_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_23_source_20_source_empty_data;
  reg _stream_matmul_23_source_21_idle;
  reg [33-1:0] _stream_matmul_23_source_21_source_count;
  reg [5-1:0] _stream_matmul_23_source_21_source_mode;
  reg [16-1:0] _stream_matmul_23_source_21_source_generator_id;
  reg [32-1:0] _stream_matmul_23_source_21_source_offset;
  reg [33-1:0] _stream_matmul_23_source_21_source_size;
  reg [32-1:0] _stream_matmul_23_source_21_source_stride;
  reg [32-1:0] _stream_matmul_23_source_21_source_offset_buf;
  reg [33-1:0] _stream_matmul_23_source_21_source_size_buf;
  reg [32-1:0] _stream_matmul_23_source_21_source_stride_buf;
  reg [8-1:0] _stream_matmul_23_source_21_source_sel;
  reg [32-1:0] _stream_matmul_23_source_21_source_ram_raddr;
  reg _stream_matmul_23_source_21_source_ram_renable;
  wire [16-1:0] _stream_matmul_23_source_21_source_ram_rdata;
  reg _stream_matmul_23_source_21_source_fifo_deq;
  wire [16-1:0] _stream_matmul_23_source_21_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_23_source_21_source_empty_data;
  wire signed [64-1:0] add_tree_2_var0_data;
  wire signed [64-1:0] _cast_src_45;
  assign _cast_src_45 = add_tree_2_var0_data;
  wire signed [64-1:0] _cast_data_45;
  assign _cast_data_45 = _cast_src_45;
  wire signed [64-1:0] add_tree_2_sum_data;
  assign add_tree_2_sum_data = _cast_data_45;
  reg [33-1:0] _stream_matmul_23_sink_26_sink_count;
  reg [5-1:0] _stream_matmul_23_sink_26_sink_mode;
  reg [16-1:0] _stream_matmul_23_sink_26_sink_generator_id;
  reg [32-1:0] _stream_matmul_23_sink_26_sink_offset;
  reg [33-1:0] _stream_matmul_23_sink_26_sink_size;
  reg [32-1:0] _stream_matmul_23_sink_26_sink_stride;
  reg [32-1:0] _stream_matmul_23_sink_26_sink_offset_buf;
  reg [33-1:0] _stream_matmul_23_sink_26_sink_size_buf;
  reg [32-1:0] _stream_matmul_23_sink_26_sink_stride_buf;
  reg [8-1:0] _stream_matmul_23_sink_26_sink_sel;
  reg [32-1:0] _stream_matmul_23_sink_26_sink_waddr;
  reg _stream_matmul_23_sink_26_sink_wenable;
  reg [16-1:0] _stream_matmul_23_sink_26_sink_wdata;
  reg _stream_matmul_23_sink_26_sink_fifo_enq;
  reg [16-1:0] _stream_matmul_23_sink_26_sink_fifo_wdata;
  reg [16-1:0] _stream_matmul_23_sink_26_sink_immediate;
  reg [33-1:0] _stream_matmul_23_sink_27_sink_count;
  reg [5-1:0] _stream_matmul_23_sink_27_sink_mode;
  reg [16-1:0] _stream_matmul_23_sink_27_sink_generator_id;
  reg [32-1:0] _stream_matmul_23_sink_27_sink_offset;
  reg [33-1:0] _stream_matmul_23_sink_27_sink_size;
  reg [32-1:0] _stream_matmul_23_sink_27_sink_stride;
  reg [32-1:0] _stream_matmul_23_sink_27_sink_offset_buf;
  reg [33-1:0] _stream_matmul_23_sink_27_sink_size_buf;
  reg [32-1:0] _stream_matmul_23_sink_27_sink_stride_buf;
  reg [8-1:0] _stream_matmul_23_sink_27_sink_sel;
  reg [32-1:0] _stream_matmul_23_sink_27_sink_waddr;
  reg _stream_matmul_23_sink_27_sink_wenable;
  reg [1-1:0] _stream_matmul_23_sink_27_sink_wdata;
  reg _stream_matmul_23_sink_27_sink_fifo_enq;
  reg [1-1:0] _stream_matmul_23_sink_27_sink_fifo_wdata;
  reg [1-1:0] _stream_matmul_23_sink_27_sink_immediate;
  reg _stream_matmul_33_stream_ivalid;
  wire _stream_matmul_33_stream_oready;
  wire _stream_matmul_33_stream_internal_oready;
  assign _stream_matmul_33_stream_oready = _stream_matmul_33_stream_internal_oready;
  reg [32-1:0] _stream_matmul_33_fsm;
  localparam _stream_matmul_33_fsm_init = 0;
  wire _stream_matmul_33_run_flag;
  reg _stream_matmul_33_source_start;
  wire _stream_matmul_33_source_stop;
  reg _stream_matmul_33_source_busy;
  wire _stream_matmul_33_sink_start;
  wire _stream_matmul_33_sink_stop;
  wire _stream_matmul_33_sink_busy;
  wire _stream_matmul_33_busy;
  reg _stream_matmul_33_busy_reg;
  wire _stream_matmul_33_is_root;
  assign _stream_matmul_33_is_root = 1;
  reg [9-1:0] _stream_matmul_33_parameter_0_next_parameter_data;
  reg [1-1:0] _stream_matmul_33_parameter_1_next_parameter_data;
  reg [1-1:0] _stream_matmul_33_parameter_2_next_parameter_data;
  reg [1-1:0] _stream_matmul_33_parameter_3_next_parameter_data;
  reg [2-1:0] _stream_matmul_33_parameter_4_next_parameter_data;
  reg [1-1:0] _stream_matmul_33_parameter_6_next_parameter_data;
  reg _stream_matmul_33_source_7_idle;
  reg [33-1:0] _stream_matmul_33_source_7_source_count;
  reg [5-1:0] _stream_matmul_33_source_7_source_mode;
  reg [16-1:0] _stream_matmul_33_source_7_source_generator_id;
  reg [32-1:0] _stream_matmul_33_source_7_source_offset;
  reg [33-1:0] _stream_matmul_33_source_7_source_size;
  reg [32-1:0] _stream_matmul_33_source_7_source_stride;
  reg [32-1:0] _stream_matmul_33_source_7_source_offset_buf;
  reg [33-1:0] _stream_matmul_33_source_7_source_size_buf;
  reg [32-1:0] _stream_matmul_33_source_7_source_stride_buf;
  reg [8-1:0] _stream_matmul_33_source_7_source_sel;
  reg [32-1:0] _stream_matmul_33_source_7_source_ram_raddr;
  reg _stream_matmul_33_source_7_source_ram_renable;
  wire [32-1:0] _stream_matmul_33_source_7_source_ram_rdata;
  reg _stream_matmul_33_source_7_source_fifo_deq;
  wire [32-1:0] _stream_matmul_33_source_7_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_33_source_7_source_empty_data;
  reg [1-1:0] _stream_matmul_33_parameter_8_next_parameter_data;
  reg _stream_matmul_33_source_9_idle;
  reg [33-1:0] _stream_matmul_33_source_9_source_count;
  reg [5-1:0] _stream_matmul_33_source_9_source_mode;
  reg [16-1:0] _stream_matmul_33_source_9_source_generator_id;
  reg [32-1:0] _stream_matmul_33_source_9_source_offset;
  reg [33-1:0] _stream_matmul_33_source_9_source_size;
  reg [32-1:0] _stream_matmul_33_source_9_source_stride;
  reg [32-1:0] _stream_matmul_33_source_9_source_offset_buf;
  reg [33-1:0] _stream_matmul_33_source_9_source_size_buf;
  reg [32-1:0] _stream_matmul_33_source_9_source_stride_buf;
  reg [8-1:0] _stream_matmul_33_source_9_source_sel;
  reg [32-1:0] _stream_matmul_33_source_9_source_ram_raddr;
  reg _stream_matmul_33_source_9_source_ram_renable;
  wire [32-1:0] _stream_matmul_33_source_9_source_ram_rdata;
  reg _stream_matmul_33_source_9_source_fifo_deq;
  wire [32-1:0] _stream_matmul_33_source_9_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_33_source_9_source_empty_data;
  reg [1-1:0] _stream_matmul_33_parameter_10_next_parameter_data;
  reg _stream_matmul_33_source_11_idle;
  reg [33-1:0] _stream_matmul_33_source_11_source_count;
  reg [5-1:0] _stream_matmul_33_source_11_source_mode;
  reg [16-1:0] _stream_matmul_33_source_11_source_generator_id;
  reg [32-1:0] _stream_matmul_33_source_11_source_offset;
  reg [33-1:0] _stream_matmul_33_source_11_source_size;
  reg [32-1:0] _stream_matmul_33_source_11_source_stride;
  reg [32-1:0] _stream_matmul_33_source_11_source_offset_buf;
  reg [33-1:0] _stream_matmul_33_source_11_source_size_buf;
  reg [32-1:0] _stream_matmul_33_source_11_source_stride_buf;
  reg [8-1:0] _stream_matmul_33_source_11_source_sel;
  reg [32-1:0] _stream_matmul_33_source_11_source_ram_raddr;
  reg _stream_matmul_33_source_11_source_ram_renable;
  wire [32-1:0] _stream_matmul_33_source_11_source_ram_rdata;
  reg _stream_matmul_33_source_11_source_fifo_deq;
  wire [32-1:0] _stream_matmul_33_source_11_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_33_source_11_source_empty_data;
  reg [1-1:0] _stream_matmul_33_parameter_12_next_parameter_data;
  reg _stream_matmul_33_source_13_idle;
  reg [33-1:0] _stream_matmul_33_source_13_source_count;
  reg [5-1:0] _stream_matmul_33_source_13_source_mode;
  reg [16-1:0] _stream_matmul_33_source_13_source_generator_id;
  reg [32-1:0] _stream_matmul_33_source_13_source_offset;
  reg [33-1:0] _stream_matmul_33_source_13_source_size;
  reg [32-1:0] _stream_matmul_33_source_13_source_stride;
  reg [32-1:0] _stream_matmul_33_source_13_source_offset_buf;
  reg [33-1:0] _stream_matmul_33_source_13_source_size_buf;
  reg [32-1:0] _stream_matmul_33_source_13_source_stride_buf;
  reg [8-1:0] _stream_matmul_33_source_13_source_sel;
  reg [32-1:0] _stream_matmul_33_source_13_source_ram_raddr;
  reg _stream_matmul_33_source_13_source_ram_renable;
  wire [32-1:0] _stream_matmul_33_source_13_source_ram_rdata;
  reg _stream_matmul_33_source_13_source_fifo_deq;
  wire [32-1:0] _stream_matmul_33_source_13_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_33_source_13_source_empty_data;
  reg [1-1:0] _stream_matmul_33_parameter_14_next_parameter_data;
  reg _stream_matmul_33_source_15_idle;
  reg [33-1:0] _stream_matmul_33_source_15_source_count;
  reg [5-1:0] _stream_matmul_33_source_15_source_mode;
  reg [16-1:0] _stream_matmul_33_source_15_source_generator_id;
  reg [32-1:0] _stream_matmul_33_source_15_source_offset;
  reg [33-1:0] _stream_matmul_33_source_15_source_size;
  reg [32-1:0] _stream_matmul_33_source_15_source_stride;
  reg [32-1:0] _stream_matmul_33_source_15_source_offset_buf;
  reg [33-1:0] _stream_matmul_33_source_15_source_size_buf;
  reg [32-1:0] _stream_matmul_33_source_15_source_stride_buf;
  reg [8-1:0] _stream_matmul_33_source_15_source_sel;
  reg [32-1:0] _stream_matmul_33_source_15_source_ram_raddr;
  reg _stream_matmul_33_source_15_source_ram_renable;
  wire [32-1:0] _stream_matmul_33_source_15_source_ram_rdata;
  reg _stream_matmul_33_source_15_source_fifo_deq;
  wire [32-1:0] _stream_matmul_33_source_15_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_33_source_15_source_empty_data;
  reg [1-1:0] _stream_matmul_33_parameter_16_next_parameter_data;
  reg [1-1:0] _stream_matmul_33_parameter_17_next_parameter_data;
  reg [5-1:0] _stream_matmul_33_parameter_18_next_parameter_data;
  reg [1-1:0] _stream_matmul_33_parameter_19_next_parameter_data;
  reg _stream_matmul_33_source_20_idle;
  reg [33-1:0] _stream_matmul_33_source_20_source_count;
  reg [5-1:0] _stream_matmul_33_source_20_source_mode;
  reg [16-1:0] _stream_matmul_33_source_20_source_generator_id;
  reg [32-1:0] _stream_matmul_33_source_20_source_offset;
  reg [33-1:0] _stream_matmul_33_source_20_source_size;
  reg [32-1:0] _stream_matmul_33_source_20_source_stride;
  reg [32-1:0] _stream_matmul_33_source_20_source_offset_buf;
  reg [33-1:0] _stream_matmul_33_source_20_source_size_buf;
  reg [32-1:0] _stream_matmul_33_source_20_source_stride_buf;
  reg [8-1:0] _stream_matmul_33_source_20_source_sel;
  reg [32-1:0] _stream_matmul_33_source_20_source_ram_raddr;
  reg _stream_matmul_33_source_20_source_ram_renable;
  wire [32-1:0] _stream_matmul_33_source_20_source_ram_rdata;
  reg _stream_matmul_33_source_20_source_fifo_deq;
  wire [32-1:0] _stream_matmul_33_source_20_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_33_source_20_source_empty_data;
  reg _stream_matmul_33_source_21_idle;
  reg [33-1:0] _stream_matmul_33_source_21_source_count;
  reg [5-1:0] _stream_matmul_33_source_21_source_mode;
  reg [16-1:0] _stream_matmul_33_source_21_source_generator_id;
  reg [32-1:0] _stream_matmul_33_source_21_source_offset;
  reg [33-1:0] _stream_matmul_33_source_21_source_size;
  reg [32-1:0] _stream_matmul_33_source_21_source_stride;
  reg [32-1:0] _stream_matmul_33_source_21_source_offset_buf;
  reg [33-1:0] _stream_matmul_33_source_21_source_size_buf;
  reg [32-1:0] _stream_matmul_33_source_21_source_stride_buf;
  reg [8-1:0] _stream_matmul_33_source_21_source_sel;
  reg [32-1:0] _stream_matmul_33_source_21_source_ram_raddr;
  reg _stream_matmul_33_source_21_source_ram_renable;
  wire [32-1:0] _stream_matmul_33_source_21_source_ram_rdata;
  reg _stream_matmul_33_source_21_source_fifo_deq;
  wire [32-1:0] _stream_matmul_33_source_21_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_33_source_21_source_empty_data;
  reg _stream_matmul_33_source_22_idle;
  reg [33-1:0] _stream_matmul_33_source_22_source_count;
  reg [5-1:0] _stream_matmul_33_source_22_source_mode;
  reg [16-1:0] _stream_matmul_33_source_22_source_generator_id;
  reg [32-1:0] _stream_matmul_33_source_22_source_offset;
  reg [33-1:0] _stream_matmul_33_source_22_source_size;
  reg [32-1:0] _stream_matmul_33_source_22_source_stride;
  reg [32-1:0] _stream_matmul_33_source_22_source_offset_buf;
  reg [33-1:0] _stream_matmul_33_source_22_source_size_buf;
  reg [32-1:0] _stream_matmul_33_source_22_source_stride_buf;
  reg [8-1:0] _stream_matmul_33_source_22_source_sel;
  reg [32-1:0] _stream_matmul_33_source_22_source_ram_raddr;
  reg _stream_matmul_33_source_22_source_ram_renable;
  wire [32-1:0] _stream_matmul_33_source_22_source_ram_rdata;
  reg _stream_matmul_33_source_22_source_fifo_deq;
  wire [32-1:0] _stream_matmul_33_source_22_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_33_source_22_source_empty_data;
  wire signed [64-1:0] add_tree_3_var0_data;
  wire signed [64-1:0] add_tree_3_var1_data;
  reg __add_tree_3_stream_ivalid_1;
  reg signed [64-1:0] __plusn_data_49;
  wire signed [64-1:0] add_tree_3_sum_data;
  assign add_tree_3_sum_data = __plusn_data_49;
  wire signed [64-1:0] add_tree_4_var0_data;
  wire signed [64-1:0] add_tree_4_var1_data;
  reg __add_tree_4_stream_ivalid_1;
  reg signed [64-1:0] __plusn_data_53;
  wire signed [64-1:0] add_tree_4_sum_data;
  assign add_tree_4_sum_data = __plusn_data_53;
  wire signed [64-1:0] acc_1_x_data;
  wire [7-1:0] acc_1_rshift_data;
  wire [32-1:0] acc_1_size_data;
  wire [1-1:0] acc_1__reduce_reset_data;
  reg __acc_1_stream_ivalid_1;
  reg __acc_1_stream_ivalid_2;
  reg __acc_1_stream_ivalid_3;
  reg __acc_1_stream_ivalid_4;
  reg __acc_1_stream_ivalid_5;
  reg [1-1:0] _greaterthan_data_25;
  reg [7-1:0] _minus_data_27;
  reg signed [64-1:0] _reduceadd_data_38;
  reg [33-1:0] _reduceadd_count_38;
  reg _reduceadd_prev_count_max_38;
  wire _reduceadd_reset_cond_38;
  assign _reduceadd_reset_cond_38 = acc_1__reduce_reset_data || _reduceadd_prev_count_max_38;
  wire [33-1:0] _reduceadd_current_count_38;
  assign _reduceadd_current_count_38 = (_reduceadd_reset_cond_38)? 0 : _reduceadd_count_38;
  wire signed [64-1:0] _reduceadd_current_data_38;
  assign _reduceadd_current_data_38 = (_reduceadd_reset_cond_38)? 1'sd0 : _reduceadd_data_38;
  reg [1-1:0] _pulse_data_40;
  reg [33-1:0] _pulse_count_40;
  reg _pulse_prev_count_max_40;
  wire _pulse_reset_cond_40;
  assign _pulse_reset_cond_40 = acc_1__reduce_reset_data || _pulse_prev_count_max_40;
  wire [33-1:0] _pulse_current_count_40;
  assign _pulse_current_count_40 = (_pulse_reset_cond_40)? 0 : _pulse_count_40;
  wire [1-1:0] _pulse_current_data_40;
  assign _pulse_current_data_40 = (_pulse_reset_cond_40)? 1'sd0 : _pulse_data_40;
  reg [7-1:0] __delay_data_1223__variable_23;
  reg signed [130-1:0] _sll_data_29;
  reg [1-1:0] __delay_data_1220_greaterthan_25;
  reg signed [64-1:0] __delay_data_1221_reduceadd_38;
  reg [7-1:0] __delay_data_1224__delay_1223__variable_23;
  reg [1-1:0] __delay_data_1227_pulse_40;
  reg signed [64-1:0] _cond_data_35;
  reg signed [64-1:0] __delay_data_1222__delay_1221_reduceadd_38;
  reg [7-1:0] __delay_data_1225__delay_1224__delay_1223__variable_23;
  reg [1-1:0] __delay_data_1228__delay_1227_pulse_40;
  reg signed [64-1:0] _plus_data_42;
  reg [7-1:0] __delay_data_1226__delay_1225__delay_1224____variable_23;
  reg [1-1:0] __delay_data_1229__delay_1228__delay_1227_pulse_40;
  reg signed [64-1:0] _sra_data_43;
  reg [1-1:0] __delay_data_1230__delay_1229__delay_1228__delay_1227_pulse_40;
  wire signed [64-1:0] acc_1_sum_data;
  assign acc_1_sum_data = _sra_data_43;
  wire [1-1:0] acc_1_valid_data;
  assign acc_1_valid_data = __delay_data_1230__delay_1229__delay_1228__delay_1227_pulse_40;
  wire signed [64-1:0] mul_rshift_round_clip_7_x_data;
  wire signed [16-1:0] mul_rshift_round_clip_7_y_data;
  wire [7-1:0] mul_rshift_round_clip_7_rshift_data;
  reg __mul_rshift_round_clip_7_stream_ivalid_1;
  reg __mul_rshift_round_clip_7_stream_ivalid_2;
  reg __mul_rshift_round_clip_7_stream_ivalid_3;
  reg __mul_rshift_round_clip_7_stream_ivalid_4;
  reg __mul_rshift_round_clip_7_stream_ivalid_5;
  reg __mul_rshift_round_clip_7_stream_ivalid_6;
  reg __mul_rshift_round_clip_7_stream_ivalid_7;
  reg __mul_rshift_round_clip_7_stream_ivalid_8;
  wire signed [80-1:0] _times_mul_odata_105;
  reg signed [80-1:0] _times_mul_odata_reg_105;
  wire signed [80-1:0] _times_data_105;
  assign _times_data_105 = _times_mul_odata_reg_105;
  wire _times_mul_update_105;
  assign _times_mul_update_105 = _mul_rshift_round_clip_7_stream_oready;

  multiplier_1
  _times_mul_105
  (
    .CLK(CLK),
    .update(_times_mul_update_105),
    .a(mul_rshift_round_clip_7_x_data),
    .b(mul_rshift_round_clip_7_y_data),
    .c(_times_mul_odata_105)
  );

  wire [7-1:0] _minus_data_108;
  assign _minus_data_108 = mul_rshift_round_clip_7_rshift_data - 2'sd1;
  wire signed [130-1:0] _sll_data_111;
  assign _sll_data_111 = 2'sd1 << _minus_data_108;
  wire [1-1:0] _eq_data_123;
  assign _eq_data_123 = mul_rshift_round_clip_7_rshift_data == 1'sd0;
  reg signed [130-1:0] __delay_data_1236_sll_111;
  reg [7-1:0] __delay_data_1240__variable_104;
  reg [1-1:0] __delay_data_1244_eq_123;
  reg signed [130-1:0] __delay_data_1237__delay_1236_sll_111;
  reg [7-1:0] __delay_data_1241__delay_1240__variable_104;
  reg [1-1:0] __delay_data_1245__delay_1244_eq_123;
  reg signed [130-1:0] __delay_data_1238__delay_1237__delay_1236_sll_111;
  reg [7-1:0] __delay_data_1242__delay_1241__delay_1240__variable_104;
  reg [1-1:0] __delay_data_1246__delay_1245__delay_1244_eq_123;
  reg signed [130-1:0] __delay_data_1239__delay_1238__delay_1237__delay_1236_sll_111;
  reg [7-1:0] __delay_data_1243__delay_1242__delay_1241____variable_104;
  reg [1-1:0] __delay_data_1247__delay_1246__delay_1245__delay_1244_eq_123;
  wire [1-1:0] _pointer_data_106;
  assign _pointer_data_106 = _times_data_105[8'sd79];
  wire signed [2-1:0] _cond_data_118;
  assign _cond_data_118 = (_pointer_data_106)? -2'sd1 : 1'sd0;
  wire signed [81-1:0] _plus_data_119;
  assign _plus_data_119 = _times_data_105 + __delay_data_1239__delay_1238__delay_1237__delay_1236_sll_111;
  wire signed [81-1:0] _plus_data_120;
  assign _plus_data_120 = _plus_data_119 + _cond_data_118;
  wire signed [80-1:0] _sra_data_121;
  assign _sra_data_121 = _plus_data_120 >>> __delay_data_1243__delay_1242__delay_1241____variable_104;
  reg signed [80-1:0] _cond_data_124;
  reg [1-1:0] _greaterthan_data_125;
  reg [1-1:0] _lessthan_data_129;
  reg [1-1:0] _greatereq_data_133;
  reg signed [80-1:0] __delay_data_1248_cond_124;
  reg signed [80-1:0] _cond_data_127;
  reg signed [80-1:0] _cond_data_131;
  reg [1-1:0] __delay_data_1249_greatereq_133;
  reg signed [16-1:0] _cond_data_135;
  wire signed [16-1:0] mul_rshift_round_clip_7_z_data;
  assign mul_rshift_round_clip_7_z_data = _cond_data_135;
  reg [33-1:0] _stream_matmul_33_sink_33_sink_count;
  reg [5-1:0] _stream_matmul_33_sink_33_sink_mode;
  reg [16-1:0] _stream_matmul_33_sink_33_sink_generator_id;
  reg [32-1:0] _stream_matmul_33_sink_33_sink_offset;
  reg [33-1:0] _stream_matmul_33_sink_33_sink_size;
  reg [32-1:0] _stream_matmul_33_sink_33_sink_stride;
  reg [32-1:0] _stream_matmul_33_sink_33_sink_offset_buf;
  reg [33-1:0] _stream_matmul_33_sink_33_sink_size_buf;
  reg [32-1:0] _stream_matmul_33_sink_33_sink_stride_buf;
  reg [8-1:0] _stream_matmul_33_sink_33_sink_sel;
  reg [32-1:0] _stream_matmul_33_sink_33_sink_waddr;
  reg _stream_matmul_33_sink_33_sink_wenable;
  reg [32-1:0] _stream_matmul_33_sink_33_sink_wdata;
  reg _stream_matmul_33_sink_33_sink_fifo_enq;
  reg [32-1:0] _stream_matmul_33_sink_33_sink_fifo_wdata;
  reg [32-1:0] _stream_matmul_33_sink_33_sink_immediate;
  reg [33-1:0] _stream_matmul_33_sink_34_sink_count;
  reg [5-1:0] _stream_matmul_33_sink_34_sink_mode;
  reg [16-1:0] _stream_matmul_33_sink_34_sink_generator_id;
  reg [32-1:0] _stream_matmul_33_sink_34_sink_offset;
  reg [33-1:0] _stream_matmul_33_sink_34_sink_size;
  reg [32-1:0] _stream_matmul_33_sink_34_sink_stride;
  reg [32-1:0] _stream_matmul_33_sink_34_sink_offset_buf;
  reg [33-1:0] _stream_matmul_33_sink_34_sink_size_buf;
  reg [32-1:0] _stream_matmul_33_sink_34_sink_stride_buf;
  reg [8-1:0] _stream_matmul_33_sink_34_sink_sel;
  reg [32-1:0] _stream_matmul_33_sink_34_sink_waddr;
  reg _stream_matmul_33_sink_34_sink_wenable;
  reg [1-1:0] _stream_matmul_33_sink_34_sink_wdata;
  reg _stream_matmul_33_sink_34_sink_fifo_enq;
  reg [1-1:0] _stream_matmul_33_sink_34_sink_fifo_wdata;
  reg [1-1:0] _stream_matmul_33_sink_34_sink_immediate;
  reg [32-1:0] main_fsm;
  localparam main_fsm_init = 0;
  reg [32-1:0] internal_state_counter;
  reg [32-1:0] conv2d_4_objaddr;
  reg [32-1:0] conv2d_4_arg_objaddr_0;
  reg [32-1:0] conv2d_4_arg_objaddr_1;
  reg [32-1:0] conv2d_4_arg_objaddr_2;
  reg [32-1:0] conv2d_4_arg_objaddr_3;
  reg [32-1:0] control_conv2d_4;
  localparam control_conv2d_4_init = 0;
  reg _control_conv2d_4_called;
  wire signed [32-1:0] conv2d_4_act_base_offset;
  reg signed [32-1:0] conv2d_4_act_base_offset_row;
  reg signed [32-1:0] conv2d_4_act_base_offset_bat;
  assign conv2d_4_act_base_offset = conv2d_4_act_base_offset_row + conv2d_4_act_base_offset_bat;
  reg signed [32-1:0] conv2d_4_filter_base_offset;
  reg [32-1:0] conv2d_4_next_stream_num_ops;
  wire signed [32-1:0] conv2d_4_out_base_offset;
  reg signed [32-1:0] conv2d_4_out_base_offset_val;
  reg signed [32-1:0] conv2d_4_out_base_offset_col;
  reg signed [32-1:0] conv2d_4_out_base_offset_row;
  reg signed [32-1:0] conv2d_4_out_base_offset_bat;
  reg signed [32-1:0] conv2d_4_out_base_offset_och;
  assign conv2d_4_out_base_offset = conv2d_4_out_base_offset_val + conv2d_4_out_base_offset_col + conv2d_4_out_base_offset_row + conv2d_4_out_base_offset_bat + conv2d_4_out_base_offset_och;
  reg conv2d_4_dma_flag_0;
  reg conv2d_4_dma_flag_1;
  reg conv2d_4_dma_flag_2;
  reg [32-1:0] conv2d_4_sync_comp_count;
  reg [32-1:0] conv2d_4_sync_out_count;
  reg [32-1:0] conv2d_4_write_count;
  reg [32-1:0] conv2d_4_next_out_write_size;
  reg [32-1:0] conv2d_4_col_count;
  reg [32-1:0] conv2d_4_row_count;
  reg [32-1:0] conv2d_4_bat_count;
  reg [32-1:0] conv2d_4_och_count;
  reg [2-1:0] conv2d_4_col_select;
  reg [2-1:0] conv2d_4_row_select;
  reg [32-1:0] conv2d_4_out_col_count;
  reg [32-1:0] conv2d_4_out_row_count;
  reg [32-1:0] conv2d_4_out_ram_select;
  reg [32-1:0] conv2d_4_prev_col_count;
  reg [32-1:0] conv2d_4_prev_row_count;
  reg [32-1:0] conv2d_4_prev_bat_count;
  reg [32-1:0] conv2d_4_prev_och_count;
  reg [2-1:0] conv2d_4_prev_row_select;
  reg [32-1:0] conv2d_4_stream_act_local_0;
  reg [32-1:0] conv2d_4_stream_act_local_1;
  reg [32-1:0] conv2d_4_stream_act_local_2;
  reg [32-1:0] conv2d_4_stream_act_local_3;
  reg [32-1:0] conv2d_4_stream_act_local_4;
  reg [32-1:0] conv2d_4_stream_act_local_5;
  reg [32-1:0] conv2d_4_stream_act_local_6;
  reg [32-1:0] conv2d_4_stream_act_local_7;
  reg [32-1:0] conv2d_4_stream_act_local_8;
  reg [32-1:0] conv2d_4_stream_out_local_val;
  reg [32-1:0] conv2d_4_stream_out_local_col;
  wire [32-1:0] conv2d_4_stream_out_local;
  assign conv2d_4_stream_out_local = conv2d_4_stream_out_local_val + conv2d_4_stream_out_local_col;
  reg [32-1:0] conv2d_4_act_page_comp_offset_0;
  reg [32-1:0] conv2d_4_act_page_comp_offset_1;
  reg [32-1:0] conv2d_4_act_page_comp_offset_2;
  reg [32-1:0] conv2d_4_act_page_dma_offset_0;
  reg [32-1:0] conv2d_4_act_page_dma_offset_1;
  reg [32-1:0] conv2d_4_act_page_dma_offset_2;
  reg [32-1:0] conv2d_4_filter_page_comp_offset;
  reg [32-1:0] conv2d_4_filter_page_dma_offset;
  reg conv2d_4_out_page;
  reg [32-1:0] conv2d_4_out_page_comp_offset;
  reg [32-1:0] conv2d_4_out_page_dma_offset;
  reg [32-1:0] conv2d_4_out_laddr_offset;
  reg conv2d_4_skip_read_filter;
  reg conv2d_4_skip_read_act;
  reg conv2d_4_skip_comp;
  reg conv2d_4_skip_write_out;
  wire [9-1:0] _dma_read_packed_high_local_size_54;
  assign _dma_read_packed_high_local_size_54 = cparam_conv2d_4_bias_num >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_55;
  assign _dma_read_packed_low_local_size_55 = cparam_conv2d_4_bias_num & { 1{ 1'd1 } };
  wire [9-1:0] _dma_read_packed_local_packed_size_56;
  assign _dma_read_packed_local_packed_size_56 = (_dma_read_packed_low_local_size_55 > 0)? _dma_read_packed_high_local_size_54 + 1 : _dma_read_packed_high_local_size_54;
  wire [32-1:0] mask_addr_shifted_57;
  assign mask_addr_shifted_57 = conv2d_4_arg_objaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_58;
  assign mask_addr_masked_58 = mask_addr_shifted_57 << 2;
  reg [32-1:0] _maxi_read_req_fsm;
  localparam _maxi_read_req_fsm_init = 0;
  reg [33-1:0] _maxi_read_cur_global_size;
  reg _maxi_read_cont;
  wire [8-1:0] pack_read_req_op_sel_59;
  wire [32-1:0] pack_read_req_local_addr_60;
  wire [32-1:0] pack_read_req_local_stride_61;
  wire [33-1:0] pack_read_req_local_size_62;
  wire [32-1:0] pack_read_req_local_blocksize_63;
  assign pack_read_req_op_sel_59 = _maxi_read_op_sel;
  assign pack_read_req_local_addr_60 = _maxi_read_local_addr;
  assign pack_read_req_local_stride_61 = _maxi_read_local_stride;
  assign pack_read_req_local_size_62 = _maxi_read_local_size;
  assign pack_read_req_local_blocksize_63 = _maxi_read_local_blocksize;
  wire [137-1:0] pack_read_req_packed_64;
  assign pack_read_req_packed_64 = { pack_read_req_op_sel_59, pack_read_req_local_addr_60, pack_read_req_local_stride_61, pack_read_req_local_size_62, pack_read_req_local_blocksize_63 };
  assign _maxi_read_req_fifo_wdata = ((_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full)? pack_read_req_packed_64 : 'hx;
  assign _maxi_read_req_fifo_enq = ((_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full)? (_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full && !_maxi_read_req_fifo_almost_full : 0;
  localparam _tmp_65 = 1;
  wire [_tmp_65-1:0] _tmp_66;
  assign _tmp_66 = !_maxi_read_req_fifo_almost_full;
  reg [_tmp_65-1:0] __tmp_66_1;
  wire [32-1:0] mask_addr_shifted_67;
  assign mask_addr_shifted_67 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_68;
  assign mask_addr_masked_68 = mask_addr_shifted_67 << 2;
  wire [32-1:0] mask_addr_shifted_69;
  assign mask_addr_shifted_69 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_70;
  assign mask_addr_masked_70 = mask_addr_shifted_69 << 2;
  wire [32-1:0] mask_addr_shifted_71;
  assign mask_addr_shifted_71 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_72;
  assign mask_addr_masked_72 = mask_addr_shifted_71 << 2;
  wire [32-1:0] mask_addr_shifted_73;
  assign mask_addr_shifted_73 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_74;
  assign mask_addr_masked_74 = mask_addr_shifted_73 << 2;
  wire [32-1:0] mask_addr_shifted_75;
  assign mask_addr_shifted_75 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_76;
  assign mask_addr_masked_76 = mask_addr_shifted_75 << 2;
  wire [32-1:0] mask_addr_shifted_77;
  assign mask_addr_shifted_77 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_78;
  assign mask_addr_masked_78 = mask_addr_shifted_77 << 2;
  reg _maxi_raddr_cond_0_1;
  reg [32-1:0] _maxi_read_data_fsm;
  localparam _maxi_read_data_fsm_init = 0;
  reg [32-1:0] write_burst_packed_fsm_0;
  localparam write_burst_packed_fsm_0_init = 0;
  reg [9-1:0] write_burst_packed_addr_79;
  reg [9-1:0] write_burst_packed_stride_80;
  reg [33-1:0] write_burst_packed_length_81;
  reg write_burst_packed_done_82;
  wire [8-1:0] write_burst_packed_ram_addr_83;
  assign write_burst_packed_ram_addr_83 = write_burst_packed_addr_79 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_84;
  assign write_burst_packed_ram_wdata_84 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id1_0_1_addr = ((write_burst_packed_fsm_0 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_83 : 'hx;
  assign ram_w16_l512_id1_0_1_wdata = ((write_burst_packed_fsm_0 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_84 : 'hx;
  assign ram_w16_l512_id1_0_1_wenable = ((write_burst_packed_fsm_0 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l512_id1_0_1_enable = ((write_burst_packed_fsm_0 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_85;
  assign write_burst_packed_ram_addr_85 = write_burst_packed_addr_79 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_86;
  assign write_burst_packed_ram_wdata_86 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id1_1_1_addr = ((write_burst_packed_fsm_0 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_85 : 'hx;
  assign ram_w16_l512_id1_1_1_wdata = ((write_burst_packed_fsm_0 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_86 : 'hx;
  assign ram_w16_l512_id1_1_1_wenable = ((write_burst_packed_fsm_0 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l512_id1_1_1_enable = ((write_burst_packed_fsm_0 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [9-1:0] _dma_read_packed_high_local_size_87;
  assign _dma_read_packed_high_local_size_87 = cparam_conv2d_4_scale_num >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_88;
  assign _dma_read_packed_low_local_size_88 = cparam_conv2d_4_scale_num & { 1{ 1'd1 } };
  wire [9-1:0] _dma_read_packed_local_packed_size_89;
  assign _dma_read_packed_local_packed_size_89 = (_dma_read_packed_low_local_size_88 > 0)? _dma_read_packed_high_local_size_87 + 1 : _dma_read_packed_high_local_size_87;
  wire [32-1:0] mask_addr_shifted_90;
  assign mask_addr_shifted_90 = conv2d_4_arg_objaddr_3 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_91;
  assign mask_addr_masked_91 = mask_addr_shifted_90 << 2;
  reg [32-1:0] write_burst_packed_fsm_1;
  localparam write_burst_packed_fsm_1_init = 0;
  reg [9-1:0] write_burst_packed_addr_92;
  reg [9-1:0] write_burst_packed_stride_93;
  reg [33-1:0] write_burst_packed_length_94;
  reg write_burst_packed_done_95;
  wire [8-1:0] write_burst_packed_ram_addr_96;
  assign write_burst_packed_ram_addr_96 = write_burst_packed_addr_92 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_97;
  assign write_burst_packed_ram_wdata_97 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id2_0_1_addr = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_96 : 'hx;
  assign ram_w16_l512_id2_0_1_wdata = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_97 : 'hx;
  assign ram_w16_l512_id2_0_1_wenable = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l512_id2_0_1_enable = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_98;
  assign write_burst_packed_ram_addr_98 = write_burst_packed_addr_92 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_99;
  assign write_burst_packed_ram_wdata_99 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id2_1_1_addr = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_98 : 'hx;
  assign ram_w16_l512_id2_1_1_wdata = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_99 : 'hx;
  assign ram_w16_l512_id2_1_1_wenable = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l512_id2_1_1_enable = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [12-1:0] _dma_write_block_high_local_size_100;
  assign _dma_write_block_high_local_size_100 = cparam_conv2d_4_filter_read_size >> 1;
  wire [1-1:0] _dma_write_block_low_local_size_101;
  assign _dma_write_block_low_local_size_101 = cparam_conv2d_4_filter_read_size & { 1{ 1'd1 } };
  wire [12-1:0] _dma_write_block_local_size_102;
  assign _dma_write_block_local_size_102 = (_dma_write_block_low_local_size_101 > 0)? _dma_write_block_high_local_size_100 + 1 : _dma_write_block_high_local_size_100;
  wire [8-1:0] _dma_read_block_high_local_blocksize_103;
  assign _dma_read_block_high_local_blocksize_103 = cparam_conv2d_4_filter_read_block >> 1;
  wire [2-1:0] _dma_read_block_low_local_blocksize_104;
  assign _dma_read_block_low_local_blocksize_104 = cparam_conv2d_4_filter_read_block & { 1{ 1'd1 } };
  wire [8-1:0] _dma_read_block_local_blocksize_105;
  assign _dma_read_block_local_blocksize_105 = (_dma_read_block_low_local_blocksize_104 > 0)? _dma_read_block_high_local_blocksize_103 + 1 : _dma_read_block_high_local_blocksize_103;
  wire [32-1:0] mask_addr_shifted_106;
  assign mask_addr_shifted_106 = conv2d_4_arg_objaddr_1 + conv2d_4_filter_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_107;
  assign mask_addr_masked_107 = mask_addr_shifted_106 << 2;
  wire write_burst_block_ram_wvalid_108;
  wire write_burst_block_ram_wquit_109;
  reg [32-1:0] write_burst_packed_fsm_2;
  localparam write_burst_packed_fsm_2_init = 0;
  reg [9-1:0] write_burst_packed_addr_110;
  reg [9-1:0] write_burst_packed_stride_111;
  reg [33-1:0] write_burst_packed_length_112;
  reg write_burst_packed_done_113;
  wire [8-1:0] write_burst_packed_ram_addr_114;
  assign write_burst_packed_ram_addr_114 = write_burst_packed_addr_110 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_115;
  assign write_burst_packed_ram_wdata_115 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id3_0_1_addr = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_108)? write_burst_packed_ram_addr_114 : 'hx;
  assign ram_w16_l512_id3_0_1_wdata = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_108)? write_burst_packed_ram_wdata_115 : 'hx;
  assign ram_w16_l512_id3_0_1_wenable = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_108)? 1'd1 : 0;
  assign ram_w16_l512_id3_0_1_enable = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_108)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_116;
  assign write_burst_packed_ram_addr_116 = write_burst_packed_addr_110 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_117;
  assign write_burst_packed_ram_wdata_117 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id3_1_1_addr = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_108)? write_burst_packed_ram_addr_116 : 'hx;
  assign ram_w16_l512_id3_1_1_wdata = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_108)? write_burst_packed_ram_wdata_117 : 'hx;
  assign ram_w16_l512_id3_1_1_wenable = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_108)? 1'd1 : 0;
  assign ram_w16_l512_id3_1_1_enable = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_108)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_118;
  wire write_burst_block_ram_wquit_119;
  reg [32-1:0] write_burst_packed_fsm_3;
  localparam write_burst_packed_fsm_3_init = 0;
  reg [9-1:0] write_burst_packed_addr_120;
  reg [9-1:0] write_burst_packed_stride_121;
  reg [33-1:0] write_burst_packed_length_122;
  reg write_burst_packed_done_123;
  wire [8-1:0] write_burst_packed_ram_addr_124;
  assign write_burst_packed_ram_addr_124 = write_burst_packed_addr_120 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_125;
  assign write_burst_packed_ram_wdata_125 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id4_0_1_addr = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_118)? write_burst_packed_ram_addr_124 : 'hx;
  assign ram_w16_l512_id4_0_1_wdata = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_118)? write_burst_packed_ram_wdata_125 : 'hx;
  assign ram_w16_l512_id4_0_1_wenable = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_118)? 1'd1 : 0;
  assign ram_w16_l512_id4_0_1_enable = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_118)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_126;
  assign write_burst_packed_ram_addr_126 = write_burst_packed_addr_120 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_127;
  assign write_burst_packed_ram_wdata_127 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id4_1_1_addr = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_118)? write_burst_packed_ram_addr_126 : 'hx;
  assign ram_w16_l512_id4_1_1_wdata = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_118)? write_burst_packed_ram_wdata_127 : 'hx;
  assign ram_w16_l512_id4_1_1_wenable = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_118)? 1'd1 : 0;
  assign ram_w16_l512_id4_1_1_enable = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_118)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_128;
  wire write_burst_block_ram_wquit_129;
  reg [32-1:0] write_burst_packed_fsm_4;
  localparam write_burst_packed_fsm_4_init = 0;
  reg [9-1:0] write_burst_packed_addr_130;
  reg [9-1:0] write_burst_packed_stride_131;
  reg [33-1:0] write_burst_packed_length_132;
  reg write_burst_packed_done_133;
  wire [8-1:0] write_burst_packed_ram_addr_134;
  assign write_burst_packed_ram_addr_134 = write_burst_packed_addr_130 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_135;
  assign write_burst_packed_ram_wdata_135 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id5_0_1_addr = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_128)? write_burst_packed_ram_addr_134 : 'hx;
  assign ram_w16_l512_id5_0_1_wdata = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_128)? write_burst_packed_ram_wdata_135 : 'hx;
  assign ram_w16_l512_id5_0_1_wenable = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_128)? 1'd1 : 0;
  assign ram_w16_l512_id5_0_1_enable = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_128)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_136;
  assign write_burst_packed_ram_addr_136 = write_burst_packed_addr_130 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_137;
  assign write_burst_packed_ram_wdata_137 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id5_1_1_addr = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_128)? write_burst_packed_ram_addr_136 : 'hx;
  assign ram_w16_l512_id5_1_1_wdata = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_128)? write_burst_packed_ram_wdata_137 : 'hx;
  assign ram_w16_l512_id5_1_1_wenable = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_128)? 1'd1 : 0;
  assign ram_w16_l512_id5_1_1_enable = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_128)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_138;
  wire write_burst_block_ram_wquit_139;
  reg [32-1:0] write_burst_packed_fsm_5;
  localparam write_burst_packed_fsm_5_init = 0;
  reg [9-1:0] write_burst_packed_addr_140;
  reg [9-1:0] write_burst_packed_stride_141;
  reg [33-1:0] write_burst_packed_length_142;
  reg write_burst_packed_done_143;
  wire [8-1:0] write_burst_packed_ram_addr_144;
  assign write_burst_packed_ram_addr_144 = write_burst_packed_addr_140 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_145;
  assign write_burst_packed_ram_wdata_145 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id6_0_1_addr = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_138)? write_burst_packed_ram_addr_144 : 'hx;
  assign ram_w16_l512_id6_0_1_wdata = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_138)? write_burst_packed_ram_wdata_145 : 'hx;
  assign ram_w16_l512_id6_0_1_wenable = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_138)? 1'd1 : 0;
  assign ram_w16_l512_id6_0_1_enable = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_138)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_146;
  assign write_burst_packed_ram_addr_146 = write_burst_packed_addr_140 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_147;
  assign write_burst_packed_ram_wdata_147 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id6_1_1_addr = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_138)? write_burst_packed_ram_addr_146 : 'hx;
  assign ram_w16_l512_id6_1_1_wdata = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_138)? write_burst_packed_ram_wdata_147 : 'hx;
  assign ram_w16_l512_id6_1_1_wenable = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_138)? 1'd1 : 0;
  assign ram_w16_l512_id6_1_1_enable = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_138)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_148;
  wire write_burst_block_ram_wquit_149;
  reg [32-1:0] write_burst_packed_fsm_6;
  localparam write_burst_packed_fsm_6_init = 0;
  reg [9-1:0] write_burst_packed_addr_150;
  reg [9-1:0] write_burst_packed_stride_151;
  reg [33-1:0] write_burst_packed_length_152;
  reg write_burst_packed_done_153;
  wire [8-1:0] write_burst_packed_ram_addr_154;
  assign write_burst_packed_ram_addr_154 = write_burst_packed_addr_150 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_155;
  assign write_burst_packed_ram_wdata_155 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id7_0_1_addr = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_148)? write_burst_packed_ram_addr_154 : 'hx;
  assign ram_w16_l512_id7_0_1_wdata = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_148)? write_burst_packed_ram_wdata_155 : 'hx;
  assign ram_w16_l512_id7_0_1_wenable = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_148)? 1'd1 : 0;
  assign ram_w16_l512_id7_0_1_enable = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_148)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_156;
  assign write_burst_packed_ram_addr_156 = write_burst_packed_addr_150 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_157;
  assign write_burst_packed_ram_wdata_157 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id7_1_1_addr = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_148)? write_burst_packed_ram_addr_156 : 'hx;
  assign ram_w16_l512_id7_1_1_wdata = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_148)? write_burst_packed_ram_wdata_157 : 'hx;
  assign ram_w16_l512_id7_1_1_wenable = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_148)? 1'd1 : 0;
  assign ram_w16_l512_id7_1_1_enable = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_148)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_158;
  wire write_burst_block_ram_wquit_159;
  reg [32-1:0] write_burst_packed_fsm_7;
  localparam write_burst_packed_fsm_7_init = 0;
  reg [9-1:0] write_burst_packed_addr_160;
  reg [9-1:0] write_burst_packed_stride_161;
  reg [33-1:0] write_burst_packed_length_162;
  reg write_burst_packed_done_163;
  wire [8-1:0] write_burst_packed_ram_addr_164;
  assign write_burst_packed_ram_addr_164 = write_burst_packed_addr_160 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_165;
  assign write_burst_packed_ram_wdata_165 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id8_0_1_addr = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_158)? write_burst_packed_ram_addr_164 : 'hx;
  assign ram_w16_l512_id8_0_1_wdata = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_158)? write_burst_packed_ram_wdata_165 : 'hx;
  assign ram_w16_l512_id8_0_1_wenable = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_158)? 1'd1 : 0;
  assign ram_w16_l512_id8_0_1_enable = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_158)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_166;
  assign write_burst_packed_ram_addr_166 = write_burst_packed_addr_160 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_167;
  assign write_burst_packed_ram_wdata_167 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id8_1_1_addr = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_158)? write_burst_packed_ram_addr_166 : 'hx;
  assign ram_w16_l512_id8_1_1_wdata = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_158)? write_burst_packed_ram_wdata_167 : 'hx;
  assign ram_w16_l512_id8_1_1_wenable = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_158)? 1'd1 : 0;
  assign ram_w16_l512_id8_1_1_enable = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_158)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_168;
  wire write_burst_block_ram_wquit_169;
  reg [32-1:0] write_burst_packed_fsm_8;
  localparam write_burst_packed_fsm_8_init = 0;
  reg [9-1:0] write_burst_packed_addr_170;
  reg [9-1:0] write_burst_packed_stride_171;
  reg [33-1:0] write_burst_packed_length_172;
  reg write_burst_packed_done_173;
  wire [8-1:0] write_burst_packed_ram_addr_174;
  assign write_burst_packed_ram_addr_174 = write_burst_packed_addr_170 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_175;
  assign write_burst_packed_ram_wdata_175 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id9_0_1_addr = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_168)? write_burst_packed_ram_addr_174 : 'hx;
  assign ram_w16_l512_id9_0_1_wdata = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_168)? write_burst_packed_ram_wdata_175 : 'hx;
  assign ram_w16_l512_id9_0_1_wenable = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_168)? 1'd1 : 0;
  assign ram_w16_l512_id9_0_1_enable = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_168)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_176;
  assign write_burst_packed_ram_addr_176 = write_burst_packed_addr_170 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_177;
  assign write_burst_packed_ram_wdata_177 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id9_1_1_addr = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_168)? write_burst_packed_ram_addr_176 : 'hx;
  assign ram_w16_l512_id9_1_1_wdata = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_168)? write_burst_packed_ram_wdata_177 : 'hx;
  assign ram_w16_l512_id9_1_1_wenable = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_168)? 1'd1 : 0;
  assign ram_w16_l512_id9_1_1_enable = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_168)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_178;
  wire write_burst_block_ram_wquit_179;
  reg [32-1:0] write_burst_packed_fsm_9;
  localparam write_burst_packed_fsm_9_init = 0;
  reg [9-1:0] write_burst_packed_addr_180;
  reg [9-1:0] write_burst_packed_stride_181;
  reg [33-1:0] write_burst_packed_length_182;
  reg write_burst_packed_done_183;
  wire [8-1:0] write_burst_packed_ram_addr_184;
  assign write_burst_packed_ram_addr_184 = write_burst_packed_addr_180 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_185;
  assign write_burst_packed_ram_wdata_185 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id10_0_1_addr = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_178)? write_burst_packed_ram_addr_184 : 'hx;
  assign ram_w16_l512_id10_0_1_wdata = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_178)? write_burst_packed_ram_wdata_185 : 'hx;
  assign ram_w16_l512_id10_0_1_wenable = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_178)? 1'd1 : 0;
  assign ram_w16_l512_id10_0_1_enable = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_178)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_186;
  assign write_burst_packed_ram_addr_186 = write_burst_packed_addr_180 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_187;
  assign write_burst_packed_ram_wdata_187 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id10_1_1_addr = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_178)? write_burst_packed_ram_addr_186 : 'hx;
  assign ram_w16_l512_id10_1_1_wdata = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_178)? write_burst_packed_ram_wdata_187 : 'hx;
  assign ram_w16_l512_id10_1_1_wenable = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_178)? 1'd1 : 0;
  assign ram_w16_l512_id10_1_1_enable = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_178)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_188;
  wire write_burst_block_ram_wquit_189;
  reg [32-1:0] write_burst_packed_fsm_10;
  localparam write_burst_packed_fsm_10_init = 0;
  reg [9-1:0] write_burst_packed_addr_190;
  reg [9-1:0] write_burst_packed_stride_191;
  reg [33-1:0] write_burst_packed_length_192;
  reg write_burst_packed_done_193;
  wire [8-1:0] write_burst_packed_ram_addr_194;
  assign write_burst_packed_ram_addr_194 = write_burst_packed_addr_190 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_195;
  assign write_burst_packed_ram_wdata_195 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id11_0_1_addr = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_188)? write_burst_packed_ram_addr_194 : 'hx;
  assign ram_w16_l512_id11_0_1_wdata = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_188)? write_burst_packed_ram_wdata_195 : 'hx;
  assign ram_w16_l512_id11_0_1_wenable = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_188)? 1'd1 : 0;
  assign ram_w16_l512_id11_0_1_enable = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_188)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_196;
  assign write_burst_packed_ram_addr_196 = write_burst_packed_addr_190 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_197;
  assign write_burst_packed_ram_wdata_197 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id11_1_1_addr = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_188)? write_burst_packed_ram_addr_196 : 'hx;
  assign ram_w16_l512_id11_1_1_wdata = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_188)? write_burst_packed_ram_wdata_197 : 'hx;
  assign ram_w16_l512_id11_1_1_wenable = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_188)? 1'd1 : 0;
  assign ram_w16_l512_id11_1_1_enable = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_188)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_11;
  localparam write_burst_block_fsm_11_init = 0;
  reg [33-1:0] write_burst_block_length_198;
  reg [32-1:0] write_burst_block_blocksize_199;
  reg write_burst_block_done_200;
  reg [32-1:0] write_burst_block_count_201;
  assign write_burst_block_ram_wvalid_108 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 1);
  assign write_burst_block_ram_wquit_109 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_118 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 2);
  assign write_burst_block_ram_wquit_119 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_128 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 3);
  assign write_burst_block_ram_wquit_129 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_138 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 4);
  assign write_burst_block_ram_wquit_139 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_148 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 5);
  assign write_burst_block_ram_wquit_149 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_158 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 6);
  assign write_burst_block_ram_wquit_159 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_168 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 7);
  assign write_burst_block_ram_wquit_169 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_178 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 8);
  assign write_burst_block_ram_wquit_179 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_188 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 9);
  assign write_burst_block_ram_wquit_189 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  wire [32-1:0] conv2d_4_mux_act_gaddr_0;
  assign conv2d_4_mux_act_gaddr_0 = (conv2d_4_row_select == 0)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_0) : 
                                    (conv2d_4_row_select == 1)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_2) : 
                                    (conv2d_4_row_select == 2)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_1) : 1'd0;
  wire [32-1:0] conv2d_4_mux_act_gaddr_1;
  assign conv2d_4_mux_act_gaddr_1 = (conv2d_4_row_select == 0)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_1) : 
                                    (conv2d_4_row_select == 1)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_0) : 
                                    (conv2d_4_row_select == 2)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_2) : 1'd0;
  wire [32-1:0] conv2d_4_mux_act_gaddr_2;
  assign conv2d_4_mux_act_gaddr_2 = (conv2d_4_row_select == 0)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_2) : 
                                    (conv2d_4_row_select == 1)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_1) : 
                                    (conv2d_4_row_select == 2)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_0) : 1'd0;
  wire conv2d_4_dma_pad_mask_0;
  assign conv2d_4_dma_pad_mask_0 = (conv2d_4_row_count + 0 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count + 0 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_dma_pad_mask_1;
  assign conv2d_4_dma_pad_mask_1 = (conv2d_4_row_count + 1 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count + 1 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_dma_pad_mask_2;
  assign conv2d_4_dma_pad_mask_2 = (conv2d_4_row_count + 2 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count + 2 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_mux_dma_pad_mask_0;
  assign conv2d_4_mux_dma_pad_mask_0 = (conv2d_4_row_select == 0)? conv2d_4_dma_pad_mask_0 : 
                                       (conv2d_4_row_select == 1)? conv2d_4_dma_pad_mask_2 : 
                                       (conv2d_4_row_select == 2)? conv2d_4_dma_pad_mask_1 : 1'd0;
  wire conv2d_4_mux_dma_pad_mask_1;
  assign conv2d_4_mux_dma_pad_mask_1 = (conv2d_4_row_select == 0)? conv2d_4_dma_pad_mask_1 : 
                                       (conv2d_4_row_select == 1)? conv2d_4_dma_pad_mask_0 : 
                                       (conv2d_4_row_select == 2)? conv2d_4_dma_pad_mask_2 : 1'd0;
  wire conv2d_4_mux_dma_pad_mask_2;
  assign conv2d_4_mux_dma_pad_mask_2 = (conv2d_4_row_select == 0)? conv2d_4_dma_pad_mask_2 : 
                                       (conv2d_4_row_select == 1)? conv2d_4_dma_pad_mask_1 : 
                                       (conv2d_4_row_select == 2)? conv2d_4_dma_pad_mask_0 : 1'd0;
  wire conv2d_4_mux_dma_flag_0;
  assign conv2d_4_mux_dma_flag_0 = (conv2d_4_prev_row_select == 0)? conv2d_4_dma_flag_0 : 
                                   (conv2d_4_prev_row_select == 1)? conv2d_4_dma_flag_2 : 
                                   (conv2d_4_prev_row_select == 2)? conv2d_4_dma_flag_1 : 1'd0;
  wire conv2d_4_mux_dma_flag_1;
  assign conv2d_4_mux_dma_flag_1 = (conv2d_4_prev_row_select == 0)? conv2d_4_dma_flag_1 : 
                                   (conv2d_4_prev_row_select == 1)? conv2d_4_dma_flag_0 : 
                                   (conv2d_4_prev_row_select == 2)? conv2d_4_dma_flag_2 : 1'd0;
  wire conv2d_4_mux_dma_flag_2;
  assign conv2d_4_mux_dma_flag_2 = (conv2d_4_prev_row_select == 0)? conv2d_4_dma_flag_2 : 
                                   (conv2d_4_prev_row_select == 1)? conv2d_4_dma_flag_1 : 
                                   (conv2d_4_prev_row_select == 2)? conv2d_4_dma_flag_0 : 1'd0;
  wire [11-1:0] _dma_write_block_high_local_size_202;
  assign _dma_write_block_high_local_size_202 = cparam_conv2d_4_act_read_size >> 1;
  wire [1-1:0] _dma_write_block_low_local_size_203;
  assign _dma_write_block_low_local_size_203 = cparam_conv2d_4_act_read_size & { 1{ 1'd1 } };
  wire [11-1:0] _dma_write_block_local_size_204;
  assign _dma_write_block_local_size_204 = (_dma_write_block_low_local_size_203 > 0)? _dma_write_block_high_local_size_202 + 1 : _dma_write_block_high_local_size_202;
  wire [8-1:0] _dma_read_block_high_local_blocksize_205;
  assign _dma_read_block_high_local_blocksize_205 = cparam_conv2d_4_act_read_block >> 1;
  wire [2-1:0] _dma_read_block_low_local_blocksize_206;
  assign _dma_read_block_low_local_blocksize_206 = cparam_conv2d_4_act_read_block & { 1{ 1'd1 } };
  wire [8-1:0] _dma_read_block_local_blocksize_207;
  assign _dma_read_block_local_blocksize_207 = (_dma_read_block_low_local_blocksize_206 > 0)? _dma_read_block_high_local_blocksize_205 + 1 : _dma_read_block_high_local_blocksize_205;
  wire [32-1:0] mask_addr_shifted_208;
  assign mask_addr_shifted_208 = conv2d_4_mux_act_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_209;
  assign mask_addr_masked_209 = mask_addr_shifted_208 << 2;
  wire write_burst_block_ram_wvalid_210;
  wire write_burst_block_ram_wquit_211;
  reg [32-1:0] write_burst_packed_fsm_12;
  localparam write_burst_packed_fsm_12_init = 0;
  reg [10-1:0] write_burst_packed_addr_212;
  reg [10-1:0] write_burst_packed_stride_213;
  reg [33-1:0] write_burst_packed_length_214;
  reg write_burst_packed_done_215;
  wire [9-1:0] write_burst_packed_ram_addr_216;
  assign write_burst_packed_ram_addr_216 = write_burst_packed_addr_212 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_217;
  assign write_burst_packed_ram_wdata_217 = _maxi_rdata_sb_0 >> 0;
  wire [9-1:0] write_burst_packed_ram_addr_218;
  assign write_burst_packed_ram_addr_218 = write_burst_packed_addr_212 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_219;
  assign write_burst_packed_ram_wdata_219 = _maxi_rdata_sb_0 >> 16;
  wire write_burst_block_ram_wvalid_220;
  wire write_burst_block_ram_wquit_221;
  reg [32-1:0] write_burst_packed_fsm_13;
  localparam write_burst_packed_fsm_13_init = 0;
  reg [10-1:0] write_burst_packed_addr_222;
  reg [10-1:0] write_burst_packed_stride_223;
  reg [33-1:0] write_burst_packed_length_224;
  reg write_burst_packed_done_225;
  wire [9-1:0] write_burst_packed_ram_addr_226;
  assign write_burst_packed_ram_addr_226 = write_burst_packed_addr_222 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_227;
  assign write_burst_packed_ram_wdata_227 = _maxi_rdata_sb_0 >> 0;
  wire [9-1:0] write_burst_packed_ram_addr_228;
  assign write_burst_packed_ram_addr_228 = write_burst_packed_addr_222 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_229;
  assign write_burst_packed_ram_wdata_229 = _maxi_rdata_sb_0 >> 16;
  wire write_burst_block_ram_wvalid_230;
  wire write_burst_block_ram_wquit_231;
  reg [32-1:0] write_burst_packed_fsm_14;
  localparam write_burst_packed_fsm_14_init = 0;
  reg [10-1:0] write_burst_packed_addr_232;
  reg [10-1:0] write_burst_packed_stride_233;
  reg [33-1:0] write_burst_packed_length_234;
  reg write_burst_packed_done_235;
  wire [9-1:0] write_burst_packed_ram_addr_236;
  assign write_burst_packed_ram_addr_236 = write_burst_packed_addr_232 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_237;
  assign write_burst_packed_ram_wdata_237 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l1024_id2_0_1_addr = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_230)? write_burst_packed_ram_addr_236 : 'hx;
  assign ram_w16_l1024_id2_0_1_wdata = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_230)? write_burst_packed_ram_wdata_237 : 'hx;
  assign ram_w16_l1024_id2_0_1_wenable = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_230)? 1'd1 : 0;
  assign ram_w16_l1024_id2_0_1_enable = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_230)? 1'd1 : 0;
  wire [9-1:0] write_burst_packed_ram_addr_238;
  assign write_burst_packed_ram_addr_238 = write_burst_packed_addr_232 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_239;
  assign write_burst_packed_ram_wdata_239 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l1024_id2_1_1_addr = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_230)? write_burst_packed_ram_addr_238 : 'hx;
  assign ram_w16_l1024_id2_1_1_wdata = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_230)? write_burst_packed_ram_wdata_239 : 'hx;
  assign ram_w16_l1024_id2_1_1_wenable = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_230)? 1'd1 : 0;
  assign ram_w16_l1024_id2_1_1_enable = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_230)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_15;
  localparam write_burst_block_fsm_15_init = 0;
  reg [33-1:0] write_burst_block_length_240;
  reg [32-1:0] write_burst_block_blocksize_241;
  reg write_burst_block_done_242;
  reg [32-1:0] write_burst_block_count_243;
  assign write_burst_block_ram_wvalid_210 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_15 == 1);
  assign write_burst_block_ram_wquit_211 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1);
  assign write_burst_block_ram_wvalid_220 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_15 == 2);
  assign write_burst_block_ram_wquit_221 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1);
  assign write_burst_block_ram_wvalid_230 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_15 == 3);
  assign write_burst_block_ram_wquit_231 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1);
  wire [11-1:0] _dma_write_block_high_local_size_244;
  assign _dma_write_block_high_local_size_244 = cparam_conv2d_4_act_read_size >> 1;
  wire [1-1:0] _dma_write_block_low_local_size_245;
  assign _dma_write_block_low_local_size_245 = cparam_conv2d_4_act_read_size & { 1{ 1'd1 } };
  wire [11-1:0] _dma_write_block_local_size_246;
  assign _dma_write_block_local_size_246 = (_dma_write_block_low_local_size_245 > 0)? _dma_write_block_high_local_size_244 + 1 : _dma_write_block_high_local_size_244;
  wire [8-1:0] _dma_read_block_high_local_blocksize_247;
  assign _dma_read_block_high_local_blocksize_247 = cparam_conv2d_4_act_read_block >> 1;
  wire [2-1:0] _dma_read_block_low_local_blocksize_248;
  assign _dma_read_block_low_local_blocksize_248 = cparam_conv2d_4_act_read_block & { 1{ 1'd1 } };
  wire [8-1:0] _dma_read_block_local_blocksize_249;
  assign _dma_read_block_local_blocksize_249 = (_dma_read_block_low_local_blocksize_248 > 0)? _dma_read_block_high_local_blocksize_247 + 1 : _dma_read_block_high_local_blocksize_247;
  wire [32-1:0] mask_addr_shifted_250;
  assign mask_addr_shifted_250 = conv2d_4_mux_act_gaddr_1 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_251;
  assign mask_addr_masked_251 = mask_addr_shifted_250 << 2;
  wire write_burst_block_ram_wvalid_252;
  wire write_burst_block_ram_wquit_253;
  reg [32-1:0] write_burst_packed_fsm_16;
  localparam write_burst_packed_fsm_16_init = 0;
  reg [10-1:0] write_burst_packed_addr_254;
  reg [10-1:0] write_burst_packed_stride_255;
  reg [33-1:0] write_burst_packed_length_256;
  reg write_burst_packed_done_257;
  wire [9-1:0] write_burst_packed_ram_addr_258;
  assign write_burst_packed_ram_addr_258 = write_burst_packed_addr_254 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_259;
  assign write_burst_packed_ram_wdata_259 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l1024_id3_0_1_addr = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_252)? write_burst_packed_ram_addr_258 : 'hx;
  assign ram_w16_l1024_id3_0_1_wdata = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_252)? write_burst_packed_ram_wdata_259 : 'hx;
  assign ram_w16_l1024_id3_0_1_wenable = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_252)? 1'd1 : 0;
  assign ram_w16_l1024_id3_0_1_enable = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_252)? 1'd1 : 0;
  wire [9-1:0] write_burst_packed_ram_addr_260;
  assign write_burst_packed_ram_addr_260 = write_burst_packed_addr_254 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_261;
  assign write_burst_packed_ram_wdata_261 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l1024_id3_1_1_addr = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_252)? write_burst_packed_ram_addr_260 : 'hx;
  assign ram_w16_l1024_id3_1_1_wdata = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_252)? write_burst_packed_ram_wdata_261 : 'hx;
  assign ram_w16_l1024_id3_1_1_wenable = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_252)? 1'd1 : 0;
  assign ram_w16_l1024_id3_1_1_enable = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_252)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_262;
  wire write_burst_block_ram_wquit_263;
  reg [32-1:0] write_burst_packed_fsm_17;
  localparam write_burst_packed_fsm_17_init = 0;
  reg [10-1:0] write_burst_packed_addr_264;
  reg [10-1:0] write_burst_packed_stride_265;
  reg [33-1:0] write_burst_packed_length_266;
  reg write_burst_packed_done_267;
  wire [9-1:0] write_burst_packed_ram_addr_268;
  assign write_burst_packed_ram_addr_268 = write_burst_packed_addr_264 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_269;
  assign write_burst_packed_ram_wdata_269 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l1024_id4_0_1_addr = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_262)? write_burst_packed_ram_addr_268 : 'hx;
  assign ram_w16_l1024_id4_0_1_wdata = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_262)? write_burst_packed_ram_wdata_269 : 'hx;
  assign ram_w16_l1024_id4_0_1_wenable = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_262)? 1'd1 : 0;
  assign ram_w16_l1024_id4_0_1_enable = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_262)? 1'd1 : 0;
  wire [9-1:0] write_burst_packed_ram_addr_270;
  assign write_burst_packed_ram_addr_270 = write_burst_packed_addr_264 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_271;
  assign write_burst_packed_ram_wdata_271 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l1024_id4_1_1_addr = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_262)? write_burst_packed_ram_addr_270 : 'hx;
  assign ram_w16_l1024_id4_1_1_wdata = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_262)? write_burst_packed_ram_wdata_271 : 'hx;
  assign ram_w16_l1024_id4_1_1_wenable = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_262)? 1'd1 : 0;
  assign ram_w16_l1024_id4_1_1_enable = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_262)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_272;
  wire write_burst_block_ram_wquit_273;
  reg [32-1:0] write_burst_packed_fsm_18;
  localparam write_burst_packed_fsm_18_init = 0;
  reg [10-1:0] write_burst_packed_addr_274;
  reg [10-1:0] write_burst_packed_stride_275;
  reg [33-1:0] write_burst_packed_length_276;
  reg write_burst_packed_done_277;
  wire [9-1:0] write_burst_packed_ram_addr_278;
  assign write_burst_packed_ram_addr_278 = write_burst_packed_addr_274 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_279;
  assign write_burst_packed_ram_wdata_279 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l1024_id5_0_1_addr = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_272)? write_burst_packed_ram_addr_278 : 'hx;
  assign ram_w16_l1024_id5_0_1_wdata = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_272)? write_burst_packed_ram_wdata_279 : 'hx;
  assign ram_w16_l1024_id5_0_1_wenable = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_272)? 1'd1 : 0;
  assign ram_w16_l1024_id5_0_1_enable = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_272)? 1'd1 : 0;
  wire [9-1:0] write_burst_packed_ram_addr_280;
  assign write_burst_packed_ram_addr_280 = write_burst_packed_addr_274 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_281;
  assign write_burst_packed_ram_wdata_281 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l1024_id5_1_1_addr = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_272)? write_burst_packed_ram_addr_280 : 'hx;
  assign ram_w16_l1024_id5_1_1_wdata = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_272)? write_burst_packed_ram_wdata_281 : 'hx;
  assign ram_w16_l1024_id5_1_1_wenable = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_272)? 1'd1 : 0;
  assign ram_w16_l1024_id5_1_1_enable = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_272)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_19;
  localparam write_burst_block_fsm_19_init = 0;
  reg [33-1:0] write_burst_block_length_282;
  reg [32-1:0] write_burst_block_blocksize_283;
  reg write_burst_block_done_284;
  reg [32-1:0] write_burst_block_count_285;
  assign write_burst_block_ram_wvalid_252 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_19 == 1);
  assign write_burst_block_ram_wquit_253 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1);
  assign write_burst_block_ram_wvalid_262 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_19 == 2);
  assign write_burst_block_ram_wquit_263 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1);
  assign write_burst_block_ram_wvalid_272 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_19 == 3);
  assign write_burst_block_ram_wquit_273 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1);
  wire [11-1:0] _dma_write_block_high_local_size_286;
  assign _dma_write_block_high_local_size_286 = cparam_conv2d_4_act_read_size >> 1;
  wire [1-1:0] _dma_write_block_low_local_size_287;
  assign _dma_write_block_low_local_size_287 = cparam_conv2d_4_act_read_size & { 1{ 1'd1 } };
  wire [11-1:0] _dma_write_block_local_size_288;
  assign _dma_write_block_local_size_288 = (_dma_write_block_low_local_size_287 > 0)? _dma_write_block_high_local_size_286 + 1 : _dma_write_block_high_local_size_286;
  wire [8-1:0] _dma_read_block_high_local_blocksize_289;
  assign _dma_read_block_high_local_blocksize_289 = cparam_conv2d_4_act_read_block >> 1;
  wire [2-1:0] _dma_read_block_low_local_blocksize_290;
  assign _dma_read_block_low_local_blocksize_290 = cparam_conv2d_4_act_read_block & { 1{ 1'd1 } };
  wire [8-1:0] _dma_read_block_local_blocksize_291;
  assign _dma_read_block_local_blocksize_291 = (_dma_read_block_low_local_blocksize_290 > 0)? _dma_read_block_high_local_blocksize_289 + 1 : _dma_read_block_high_local_blocksize_289;
  wire [32-1:0] mask_addr_shifted_292;
  assign mask_addr_shifted_292 = conv2d_4_mux_act_gaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_293;
  assign mask_addr_masked_293 = mask_addr_shifted_292 << 2;
  wire write_burst_block_ram_wvalid_294;
  wire write_burst_block_ram_wquit_295;
  reg [32-1:0] write_burst_packed_fsm_20;
  localparam write_burst_packed_fsm_20_init = 0;
  reg [10-1:0] write_burst_packed_addr_296;
  reg [10-1:0] write_burst_packed_stride_297;
  reg [33-1:0] write_burst_packed_length_298;
  reg write_burst_packed_done_299;
  wire [9-1:0] write_burst_packed_ram_addr_300;
  assign write_burst_packed_ram_addr_300 = write_burst_packed_addr_296 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_301;
  assign write_burst_packed_ram_wdata_301 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l1024_id6_0_1_addr = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_294)? write_burst_packed_ram_addr_300 : 'hx;
  assign ram_w16_l1024_id6_0_1_wdata = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_294)? write_burst_packed_ram_wdata_301 : 'hx;
  assign ram_w16_l1024_id6_0_1_wenable = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_294)? 1'd1 : 0;
  assign ram_w16_l1024_id6_0_1_enable = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_294)? 1'd1 : 0;
  wire [9-1:0] write_burst_packed_ram_addr_302;
  assign write_burst_packed_ram_addr_302 = write_burst_packed_addr_296 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_303;
  assign write_burst_packed_ram_wdata_303 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l1024_id6_1_1_addr = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_294)? write_burst_packed_ram_addr_302 : 'hx;
  assign ram_w16_l1024_id6_1_1_wdata = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_294)? write_burst_packed_ram_wdata_303 : 'hx;
  assign ram_w16_l1024_id6_1_1_wenable = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_294)? 1'd1 : 0;
  assign ram_w16_l1024_id6_1_1_enable = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_294)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_304;
  wire write_burst_block_ram_wquit_305;
  reg [32-1:0] write_burst_packed_fsm_21;
  localparam write_burst_packed_fsm_21_init = 0;
  reg [10-1:0] write_burst_packed_addr_306;
  reg [10-1:0] write_burst_packed_stride_307;
  reg [33-1:0] write_burst_packed_length_308;
  reg write_burst_packed_done_309;
  wire [9-1:0] write_burst_packed_ram_addr_310;
  assign write_burst_packed_ram_addr_310 = write_burst_packed_addr_306 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_311;
  assign write_burst_packed_ram_wdata_311 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l1024_id7_0_1_addr = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_304)? write_burst_packed_ram_addr_310 : 'hx;
  assign ram_w16_l1024_id7_0_1_wdata = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_304)? write_burst_packed_ram_wdata_311 : 'hx;
  assign ram_w16_l1024_id7_0_1_wenable = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_304)? 1'd1 : 0;
  assign ram_w16_l1024_id7_0_1_enable = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_304)? 1'd1 : 0;
  wire [9-1:0] write_burst_packed_ram_addr_312;
  assign write_burst_packed_ram_addr_312 = write_burst_packed_addr_306 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_313;
  assign write_burst_packed_ram_wdata_313 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l1024_id7_1_1_addr = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_304)? write_burst_packed_ram_addr_312 : 'hx;
  assign ram_w16_l1024_id7_1_1_wdata = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_304)? write_burst_packed_ram_wdata_313 : 'hx;
  assign ram_w16_l1024_id7_1_1_wenable = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_304)? 1'd1 : 0;
  assign ram_w16_l1024_id7_1_1_enable = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_304)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_314;
  wire write_burst_block_ram_wquit_315;
  reg [32-1:0] write_burst_packed_fsm_22;
  localparam write_burst_packed_fsm_22_init = 0;
  reg [10-1:0] write_burst_packed_addr_316;
  reg [10-1:0] write_burst_packed_stride_317;
  reg [33-1:0] write_burst_packed_length_318;
  reg write_burst_packed_done_319;
  wire [9-1:0] write_burst_packed_ram_addr_320;
  assign write_burst_packed_ram_addr_320 = write_burst_packed_addr_316 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_321;
  assign write_burst_packed_ram_wdata_321 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l1024_id8_0_1_addr = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_314)? write_burst_packed_ram_addr_320 : 'hx;
  assign ram_w16_l1024_id8_0_1_wdata = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_314)? write_burst_packed_ram_wdata_321 : 'hx;
  assign ram_w16_l1024_id8_0_1_wenable = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_314)? 1'd1 : 0;
  assign ram_w16_l1024_id8_0_1_enable = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_314)? 1'd1 : 0;
  wire [9-1:0] write_burst_packed_ram_addr_322;
  assign write_burst_packed_ram_addr_322 = write_burst_packed_addr_316 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_323;
  assign write_burst_packed_ram_wdata_323 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l1024_id8_1_1_addr = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_314)? write_burst_packed_ram_addr_322 : 'hx;
  assign ram_w16_l1024_id8_1_1_wdata = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_314)? write_burst_packed_ram_wdata_323 : 'hx;
  assign ram_w16_l1024_id8_1_1_wenable = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_314)? 1'd1 : 0;
  assign ram_w16_l1024_id8_1_1_enable = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_314)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_23;
  localparam write_burst_block_fsm_23_init = 0;
  reg [33-1:0] write_burst_block_length_324;
  reg [32-1:0] write_burst_block_blocksize_325;
  reg write_burst_block_done_326;
  reg [32-1:0] write_burst_block_count_327;
  assign write_burst_block_ram_wvalid_294 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_23 == 1);
  assign write_burst_block_ram_wquit_295 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1);
  assign write_burst_block_ram_wvalid_304 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_23 == 2);
  assign write_burst_block_ram_wquit_305 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1);
  assign write_burst_block_ram_wvalid_314 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_23 == 3);
  assign write_burst_block_ram_wquit_315 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1);
  reg [32-1:0] conv2d_4_comp_fsm;
  localparam conv2d_4_comp_fsm_init = 0;
  reg [32-1:0] conv2d_4_filter_page_comp_offset_buf;
  reg [32-1:0] conv2d_4_act_page_comp_offset_buf_0;
  reg [32-1:0] conv2d_4_act_page_comp_offset_buf_1;
  reg [32-1:0] conv2d_4_act_page_comp_offset_buf_2;
  reg [32-1:0] conv2d_4_out_page_comp_offset_buf;
  reg [32-1:0] conv2d_4_row_count_buf;
  reg [2-1:0] conv2d_4_row_select_buf;
  reg [32-1:0] conv2d_4_och_count_buf;
  wire conv2d_4_stream_pad_mask_0_0;
  assign conv2d_4_stream_pad_mask_0_0 = (conv2d_4_col_count + 0 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 0 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 0 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 0 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_0_1;
  assign conv2d_4_stream_pad_mask_0_1 = (conv2d_4_col_count + 1 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 1 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 0 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 0 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_0_2;
  assign conv2d_4_stream_pad_mask_0_2 = (conv2d_4_col_count + 2 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 2 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 0 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 0 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_1_0;
  assign conv2d_4_stream_pad_mask_1_0 = (conv2d_4_col_count + 0 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 0 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 1 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 1 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_1_1;
  assign conv2d_4_stream_pad_mask_1_1 = (conv2d_4_col_count + 1 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 1 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 1 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 1 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_1_2;
  assign conv2d_4_stream_pad_mask_1_2 = (conv2d_4_col_count + 2 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 2 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 1 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 1 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_2_0;
  assign conv2d_4_stream_pad_mask_2_0 = (conv2d_4_col_count + 0 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 0 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 2 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 2 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_2_1;
  assign conv2d_4_stream_pad_mask_2_1 = (conv2d_4_col_count + 1 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 1 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 2 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 2 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_2_2;
  assign conv2d_4_stream_pad_mask_2_2 = (conv2d_4_col_count + 2 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 2 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 2 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 2 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  reg [9-1:0] conv2d_4_stream_pad_masks;
  wire [8-1:0] stream_conv2d_4_parameter_0_data;
  wire [2-1:0] stream_conv2d_4_parameter_1_data;
  wire [2-1:0] stream_conv2d_4_parameter_2_data;
  wire [9-1:0] stream_conv2d_4_parameter_3_data;
  wire [1-1:0] stream_conv2d_4_parameter_4_data;
  wire [1-1:0] stream_conv2d_4__reduce_reset_data;
  wire [1-1:0] stream_conv2d_4_parameter_6_data;
  wire [16-1:0] stream_conv2d_4_source_7_data;
  wire [1-1:0] stream_conv2d_4_parameter_8_data;
  wire [16-1:0] stream_conv2d_4_source_9_data;
  wire [1-1:0] stream_conv2d_4_parameter_10_data;
  wire [16-1:0] stream_conv2d_4_source_11_data;
  wire [1-1:0] stream_conv2d_4_parameter_12_data;
  wire [16-1:0] stream_conv2d_4_source_13_data;
  wire [1-1:0] stream_conv2d_4_parameter_14_data;
  wire [16-1:0] stream_conv2d_4_source_15_data;
  wire [1-1:0] stream_conv2d_4_parameter_16_data;
  wire [1-1:0] stream_conv2d_4_parameter_17_data;
  wire [1-1:0] stream_conv2d_4_parameter_18_data;
  wire [1-1:0] stream_conv2d_4_parameter_19_data;
  wire [16-1:0] stream_conv2d_4_source_20_data;
  wire [16-1:0] stream_conv2d_4_source_21_data;
  wire [16-1:0] stream_conv2d_4_source_22_data;
  wire [16-1:0] stream_conv2d_4_source_23_data;
  wire [16-1:0] stream_conv2d_4_source_24_data;
  wire [16-1:0] stream_conv2d_4_source_25_data;
  wire [16-1:0] stream_conv2d_4_source_26_data;
  wire [16-1:0] stream_conv2d_4_source_27_data;
  wire [16-1:0] stream_conv2d_4_source_28_data;
  wire [16-1:0] stream_conv2d_4_source_29_data;
  wire [16-1:0] stream_conv2d_4_source_30_data;
  wire [16-1:0] stream_conv2d_4_source_31_data;
  wire [16-1:0] stream_conv2d_4_source_32_data;
  wire [16-1:0] stream_conv2d_4_source_33_data;
  wire [16-1:0] stream_conv2d_4_source_34_data;
  wire [16-1:0] stream_conv2d_4_source_35_data;
  wire [16-1:0] stream_conv2d_4_source_36_data;
  wire [16-1:0] stream_conv2d_4_source_37_data;
  reg __stream_conv2d_4_stream_ivalid_1;
  reg __stream_conv2d_4_stream_ivalid_2;
  reg __stream_conv2d_4_stream_ivalid_3;
  reg __stream_conv2d_4_stream_ivalid_4;
  reg __stream_conv2d_4_stream_ivalid_5;
  reg __stream_conv2d_4_stream_ivalid_6;
  reg __stream_conv2d_4_stream_ivalid_7;
  reg __stream_conv2d_4_stream_ivalid_8;
  reg __stream_conv2d_4_stream_ivalid_9;
  reg __stream_conv2d_4_stream_ivalid_10;
  reg __stream_conv2d_4_stream_ivalid_11;
  reg __stream_conv2d_4_stream_ivalid_12;
  reg __stream_conv2d_4_stream_ivalid_13;
  reg __stream_conv2d_4_stream_ivalid_14;
  reg __stream_conv2d_4_stream_ivalid_15;
  reg __stream_conv2d_4_stream_ivalid_16;
  reg __stream_conv2d_4_stream_ivalid_17;
  reg __stream_conv2d_4_stream_ivalid_18;
  reg __stream_conv2d_4_stream_ivalid_19;
  reg __stream_conv2d_4_stream_ivalid_20;
  reg __stream_conv2d_4_stream_ivalid_21;
  reg __stream_conv2d_4_stream_ivalid_22;
  reg __stream_conv2d_4_stream_ivalid_23;
  reg __stream_conv2d_4_stream_ivalid_24;
  reg __stream_conv2d_4_stream_ivalid_25;
  reg __stream_conv2d_4_stream_ivalid_26;
  reg __stream_conv2d_4_stream_ivalid_27;
  reg __stream_conv2d_4_stream_ivalid_28;
  reg __stream_conv2d_4_stream_ivalid_29;
  reg __stream_conv2d_4_stream_ivalid_30;
  reg __stream_conv2d_4_stream_ivalid_31;
  wire [16-1:0] _slice_data_358;
  assign _slice_data_358 = stream_conv2d_4_source_7_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_359;
  assign _reinterpretcast_src_359 = _slice_data_358;
  wire signed [16-1:0] _reinterpretcast_data_359;
  assign _reinterpretcast_data_359 = _reinterpretcast_src_359;
  wire signed [16-1:0] _cond_data_360;
  assign _cond_data_360 = (stream_conv2d_4_parameter_6_data)? _reinterpretcast_data_359 : _reinterpretcast_data_359;
  wire [16-1:0] _slice_data_365;
  assign _slice_data_365 = stream_conv2d_4_source_9_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_366;
  assign _reinterpretcast_src_366 = _slice_data_365;
  wire signed [16-1:0] _reinterpretcast_data_366;
  assign _reinterpretcast_data_366 = _reinterpretcast_src_366;
  wire signed [16-1:0] _cond_data_367;
  assign _cond_data_367 = (stream_conv2d_4_parameter_8_data)? _reinterpretcast_data_366 : _reinterpretcast_data_366;
  wire [16-1:0] _slice_data_372;
  assign _slice_data_372 = stream_conv2d_4_source_11_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_373;
  assign _reinterpretcast_src_373 = _slice_data_372;
  wire [16-1:0] _reinterpretcast_data_373;
  assign _reinterpretcast_data_373 = _reinterpretcast_src_373;
  wire [16-1:0] _cond_data_374;
  assign _cond_data_374 = (stream_conv2d_4_parameter_10_data)? _reinterpretcast_data_373 : _reinterpretcast_data_373;
  wire [16-1:0] _slice_data_379;
  assign _slice_data_379 = stream_conv2d_4_source_13_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_380;
  assign _reinterpretcast_src_380 = _slice_data_379;
  wire [16-1:0] _reinterpretcast_data_380;
  assign _reinterpretcast_data_380 = _reinterpretcast_src_380;
  wire [16-1:0] _cond_data_381;
  assign _cond_data_381 = (stream_conv2d_4_parameter_12_data)? _reinterpretcast_data_380 : _reinterpretcast_data_380;
  wire [16-1:0] _slice_data_386;
  assign _slice_data_386 = stream_conv2d_4_source_15_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_387;
  assign _reinterpretcast_src_387 = _slice_data_386;
  wire [16-1:0] _reinterpretcast_data_387;
  assign _reinterpretcast_data_387 = _reinterpretcast_src_387;
  wire [16-1:0] _cond_data_388;
  assign _cond_data_388 = (stream_conv2d_4_parameter_14_data)? _reinterpretcast_data_387 : _reinterpretcast_data_387;
  reg [1-1:0] _eq_data_402;
  reg [1-1:0] _eq_data_406;
  reg [1-1:0] _eq_data_409;
  reg [1-1:0] _eq_data_412;
  reg [1-1:0] _eq_data_416;
  reg [1-1:0] _eq_data_419;
  reg [1-1:0] _eq_data_422;
  reg [1-1:0] _eq_data_426;
  reg [1-1:0] _eq_data_429;
  reg [1-1:0] _eq_data_432;
  reg [1-1:0] _eq_data_436;
  reg [1-1:0] _eq_data_439;
  reg [1-1:0] _eq_data_442;
  reg [1-1:0] _eq_data_446;
  reg [1-1:0] _eq_data_449;
  reg [1-1:0] _eq_data_452;
  reg [1-1:0] _eq_data_456;
  reg [1-1:0] _eq_data_459;
  reg [1-1:0] _eq_data_462;
  reg [1-1:0] _eq_data_466;
  reg [1-1:0] _eq_data_469;
  reg [1-1:0] _eq_data_472;
  reg [1-1:0] _eq_data_476;
  reg [1-1:0] _eq_data_479;
  reg [1-1:0] _eq_data_482;
  reg [1-1:0] _eq_data_486;
  reg [1-1:0] _eq_data_489;
  reg [1-1:0] _eq_data_492;
  reg [1-1:0] _eq_data_496;
  reg [1-1:0] _eq_data_499;
  reg [1-1:0] _eq_data_502;
  reg [1-1:0] _eq_data_506;
  reg [1-1:0] _eq_data_509;
  reg [1-1:0] _eq_data_512;
  reg [1-1:0] _eq_data_516;
  reg [1-1:0] _eq_data_519;
  reg [1-1:0] _eq_data_522;
  reg [1-1:0] _eq_data_526;
  reg [1-1:0] _eq_data_529;
  reg [1-1:0] _eq_data_532;
  reg [1-1:0] _eq_data_536;
  reg [1-1:0] _eq_data_539;
  reg [1-1:0] _eq_data_542;
  reg [1-1:0] _eq_data_546;
  reg [1-1:0] _eq_data_549;
  reg [1-1:0] _eq_data_552;
  reg [1-1:0] _eq_data_556;
  reg [1-1:0] _eq_data_559;
  reg [1-1:0] _eq_data_562;
  reg [1-1:0] _eq_data_566;
  reg [1-1:0] _eq_data_569;
  reg [1-1:0] _eq_data_572;
  reg [1-1:0] _eq_data_576;
  reg [1-1:0] _eq_data_579;
  wire [16-1:0] _reinterpretcast_src_672;
  assign _reinterpretcast_src_672 = stream_conv2d_4_source_29_data;
  wire signed [16-1:0] _reinterpretcast_data_672;
  assign _reinterpretcast_data_672 = _reinterpretcast_src_672;
  wire [16-1:0] _reinterpretcast_src_673;
  assign _reinterpretcast_src_673 = stream_conv2d_4_source_30_data;
  wire signed [16-1:0] _reinterpretcast_data_673;
  assign _reinterpretcast_data_673 = _reinterpretcast_src_673;
  wire [16-1:0] _reinterpretcast_src_674;
  assign _reinterpretcast_src_674 = stream_conv2d_4_source_31_data;
  wire signed [16-1:0] _reinterpretcast_data_674;
  assign _reinterpretcast_data_674 = _reinterpretcast_src_674;
  wire [16-1:0] _reinterpretcast_src_675;
  assign _reinterpretcast_src_675 = stream_conv2d_4_source_32_data;
  wire signed [16-1:0] _reinterpretcast_data_675;
  assign _reinterpretcast_data_675 = _reinterpretcast_src_675;
  wire [16-1:0] _reinterpretcast_src_676;
  assign _reinterpretcast_src_676 = stream_conv2d_4_source_33_data;
  wire signed [16-1:0] _reinterpretcast_data_676;
  assign _reinterpretcast_data_676 = _reinterpretcast_src_676;
  wire [16-1:0] _reinterpretcast_src_677;
  assign _reinterpretcast_src_677 = stream_conv2d_4_source_34_data;
  wire signed [16-1:0] _reinterpretcast_data_677;
  assign _reinterpretcast_data_677 = _reinterpretcast_src_677;
  wire [16-1:0] _reinterpretcast_src_678;
  assign _reinterpretcast_src_678 = stream_conv2d_4_source_35_data;
  wire signed [16-1:0] _reinterpretcast_data_678;
  assign _reinterpretcast_data_678 = _reinterpretcast_src_678;
  wire [16-1:0] _reinterpretcast_src_679;
  assign _reinterpretcast_src_679 = stream_conv2d_4_source_36_data;
  wire signed [16-1:0] _reinterpretcast_data_679;
  assign _reinterpretcast_data_679 = _reinterpretcast_src_679;
  wire [16-1:0] _reinterpretcast_src_680;
  assign _reinterpretcast_src_680 = stream_conv2d_4_source_37_data;
  wire signed [16-1:0] _reinterpretcast_data_680;
  assign _reinterpretcast_data_680 = _reinterpretcast_src_680;
  wire [1-1:0] _pointer_data_681;
  assign _pointer_data_681 = stream_conv2d_4_parameter_3_data[1'sd0];
  wire [1-1:0] _pointer_data_683;
  assign _pointer_data_683 = stream_conv2d_4_parameter_3_data[2'sd1];
  wire [1-1:0] _pointer_data_685;
  assign _pointer_data_685 = stream_conv2d_4_parameter_3_data[3'sd2];
  wire [1-1:0] _pointer_data_687;
  assign _pointer_data_687 = stream_conv2d_4_parameter_3_data[3'sd3];
  wire [1-1:0] _pointer_data_689;
  assign _pointer_data_689 = stream_conv2d_4_parameter_3_data[4'sd4];
  wire [1-1:0] _pointer_data_691;
  assign _pointer_data_691 = stream_conv2d_4_parameter_3_data[4'sd5];
  wire [1-1:0] _pointer_data_693;
  assign _pointer_data_693 = stream_conv2d_4_parameter_3_data[4'sd6];
  wire [1-1:0] _pointer_data_695;
  assign _pointer_data_695 = stream_conv2d_4_parameter_3_data[4'sd7];
  wire [1-1:0] _pointer_data_697;
  assign _pointer_data_697 = stream_conv2d_4_parameter_3_data[5'sd8];
  reg [16-1:0] _plus_data_734;
  reg [16-1:0] _plus_data_753;
  reg [16-1:0] _plus_data_772;
  reg [16-1:0] _plus_data_791;
  reg [16-1:0] _plus_data_810;
  reg [16-1:0] _plus_data_829;
  reg [16-1:0] _plus_data_848;
  reg [16-1:0] _plus_data_867;
  reg [16-1:0] _plus_data_886;
  reg [16-1:0] _plus_data_902;
  reg [16-1:0] _plus_data_921;
  reg [16-1:0] __delay_data_1254__variable_395;
  reg [16-1:0] __delay_data_1255__variable_394;
  reg [16-1:0] __delay_data_1256__variable_393;
  reg [16-1:0] __delay_data_1257__variable_398;
  reg [16-1:0] __delay_data_1258__variable_397;
  reg [16-1:0] __delay_data_1259__variable_396;
  reg [16-1:0] __delay_data_1260__variable_401;
  reg [16-1:0] __delay_data_1261__variable_400;
  reg [16-1:0] __delay_data_1262__variable_399;
  reg [1-1:0] __delay_data_1263_pointer_681;
  reg signed [16-1:0] __delay_data_1264_reinterpretcast_672;
  reg [1-1:0] __delay_data_1265_pointer_683;
  reg signed [16-1:0] __delay_data_1266_reinterpretcast_673;
  reg [1-1:0] __delay_data_1267_pointer_685;
  reg signed [16-1:0] __delay_data_1268_reinterpretcast_674;
  reg [1-1:0] __delay_data_1269_pointer_687;
  reg signed [16-1:0] __delay_data_1270_reinterpretcast_675;
  reg [1-1:0] __delay_data_1271_pointer_689;
  reg signed [16-1:0] __delay_data_1272_reinterpretcast_676;
  reg [1-1:0] __delay_data_1273_pointer_691;
  reg signed [16-1:0] __delay_data_1274_reinterpretcast_677;
  reg [1-1:0] __delay_data_1275_pointer_693;
  reg signed [16-1:0] __delay_data_1276_reinterpretcast_678;
  reg [1-1:0] __delay_data_1277_pointer_695;
  reg signed [16-1:0] __delay_data_1278_reinterpretcast_679;
  reg [1-1:0] __delay_data_1279_pointer_697;
  reg signed [16-1:0] __delay_data_1280_reinterpretcast_680;
  reg [1-1:0] __delay_data_1281__variable_344;
  reg [8-1:0] __delay_data_1306__variable_339;
  reg signed [16-1:0] __delay_data_1319_cond_360;
  reg signed [16-1:0] __delay_data_1338_cond_367;
  wire signed [16-1:0] _cond_data_404;
  assign _cond_data_404 = (_eq_data_402)? __delay_data_1254__variable_395 : 1'sd0;
  wire signed [16-1:0] _cond_data_408;
  assign _cond_data_408 = (_eq_data_406)? __delay_data_1255__variable_394 : _cond_data_404;
  wire signed [16-1:0] _cond_data_411;
  assign _cond_data_411 = (_eq_data_409)? __delay_data_1256__variable_393 : _cond_data_408;
  wire signed [16-1:0] _cond_data_414;
  assign _cond_data_414 = (_eq_data_412)? __delay_data_1256__variable_393 : 1'sd0;
  wire signed [16-1:0] _cond_data_418;
  assign _cond_data_418 = (_eq_data_416)? __delay_data_1254__variable_395 : _cond_data_414;
  wire signed [16-1:0] _cond_data_421;
  assign _cond_data_421 = (_eq_data_419)? __delay_data_1255__variable_394 : _cond_data_418;
  wire signed [16-1:0] _cond_data_424;
  assign _cond_data_424 = (_eq_data_422)? __delay_data_1255__variable_394 : 1'sd0;
  wire signed [16-1:0] _cond_data_428;
  assign _cond_data_428 = (_eq_data_426)? __delay_data_1256__variable_393 : _cond_data_424;
  wire signed [16-1:0] _cond_data_431;
  assign _cond_data_431 = (_eq_data_429)? __delay_data_1254__variable_395 : _cond_data_428;
  wire signed [16-1:0] _cond_data_434;
  assign _cond_data_434 = (_eq_data_432)? __delay_data_1257__variable_398 : 1'sd0;
  wire signed [16-1:0] _cond_data_438;
  assign _cond_data_438 = (_eq_data_436)? __delay_data_1258__variable_397 : _cond_data_434;
  wire signed [16-1:0] _cond_data_441;
  assign _cond_data_441 = (_eq_data_439)? __delay_data_1259__variable_396 : _cond_data_438;
  wire signed [16-1:0] _cond_data_444;
  assign _cond_data_444 = (_eq_data_442)? __delay_data_1259__variable_396 : 1'sd0;
  wire signed [16-1:0] _cond_data_448;
  assign _cond_data_448 = (_eq_data_446)? __delay_data_1257__variable_398 : _cond_data_444;
  wire signed [16-1:0] _cond_data_451;
  assign _cond_data_451 = (_eq_data_449)? __delay_data_1258__variable_397 : _cond_data_448;
  wire signed [16-1:0] _cond_data_454;
  assign _cond_data_454 = (_eq_data_452)? __delay_data_1258__variable_397 : 1'sd0;
  wire signed [16-1:0] _cond_data_458;
  assign _cond_data_458 = (_eq_data_456)? __delay_data_1259__variable_396 : _cond_data_454;
  wire signed [16-1:0] _cond_data_461;
  assign _cond_data_461 = (_eq_data_459)? __delay_data_1257__variable_398 : _cond_data_458;
  wire signed [16-1:0] _cond_data_464;
  assign _cond_data_464 = (_eq_data_462)? __delay_data_1260__variable_401 : 1'sd0;
  wire signed [16-1:0] _cond_data_468;
  assign _cond_data_468 = (_eq_data_466)? __delay_data_1261__variable_400 : _cond_data_464;
  wire signed [16-1:0] _cond_data_471;
  assign _cond_data_471 = (_eq_data_469)? __delay_data_1262__variable_399 : _cond_data_468;
  wire signed [16-1:0] _cond_data_474;
  assign _cond_data_474 = (_eq_data_472)? __delay_data_1262__variable_399 : 1'sd0;
  wire signed [16-1:0] _cond_data_478;
  assign _cond_data_478 = (_eq_data_476)? __delay_data_1260__variable_401 : _cond_data_474;
  wire signed [16-1:0] _cond_data_481;
  assign _cond_data_481 = (_eq_data_479)? __delay_data_1261__variable_400 : _cond_data_478;
  wire signed [16-1:0] _cond_data_484;
  assign _cond_data_484 = (_eq_data_482)? __delay_data_1261__variable_400 : 1'sd0;
  wire signed [16-1:0] _cond_data_488;
  assign _cond_data_488 = (_eq_data_486)? __delay_data_1262__variable_399 : _cond_data_484;
  wire signed [16-1:0] _cond_data_491;
  assign _cond_data_491 = (_eq_data_489)? __delay_data_1260__variable_401 : _cond_data_488;
  wire signed [16-1:0] _cond_data_494;
  assign _cond_data_494 = (_eq_data_492)? _cond_data_471 : 1'sd0;
  wire signed [16-1:0] _cond_data_498;
  assign _cond_data_498 = (_eq_data_496)? _cond_data_441 : _cond_data_494;
  wire signed [16-1:0] _cond_data_501;
  assign _cond_data_501 = (_eq_data_499)? _cond_data_411 : _cond_data_498;
  wire signed [16-1:0] _cond_data_504;
  assign _cond_data_504 = (_eq_data_502)? _cond_data_411 : 1'sd0;
  wire signed [16-1:0] _cond_data_508;
  assign _cond_data_508 = (_eq_data_506)? _cond_data_471 : _cond_data_504;
  wire signed [16-1:0] _cond_data_511;
  assign _cond_data_511 = (_eq_data_509)? _cond_data_441 : _cond_data_508;
  wire signed [16-1:0] _cond_data_514;
  assign _cond_data_514 = (_eq_data_512)? _cond_data_441 : 1'sd0;
  wire signed [16-1:0] _cond_data_518;
  assign _cond_data_518 = (_eq_data_516)? _cond_data_411 : _cond_data_514;
  wire signed [16-1:0] _cond_data_521;
  assign _cond_data_521 = (_eq_data_519)? _cond_data_471 : _cond_data_518;
  wire signed [16-1:0] _cond_data_524;
  assign _cond_data_524 = (_eq_data_522)? _cond_data_481 : 1'sd0;
  wire signed [16-1:0] _cond_data_528;
  assign _cond_data_528 = (_eq_data_526)? _cond_data_451 : _cond_data_524;
  wire signed [16-1:0] _cond_data_531;
  assign _cond_data_531 = (_eq_data_529)? _cond_data_421 : _cond_data_528;
  wire signed [16-1:0] _cond_data_534;
  assign _cond_data_534 = (_eq_data_532)? _cond_data_421 : 1'sd0;
  wire signed [16-1:0] _cond_data_538;
  assign _cond_data_538 = (_eq_data_536)? _cond_data_481 : _cond_data_534;
  wire signed [16-1:0] _cond_data_541;
  assign _cond_data_541 = (_eq_data_539)? _cond_data_451 : _cond_data_538;
  wire signed [16-1:0] _cond_data_544;
  assign _cond_data_544 = (_eq_data_542)? _cond_data_451 : 1'sd0;
  wire signed [16-1:0] _cond_data_548;
  assign _cond_data_548 = (_eq_data_546)? _cond_data_421 : _cond_data_544;
  wire signed [16-1:0] _cond_data_551;
  assign _cond_data_551 = (_eq_data_549)? _cond_data_481 : _cond_data_548;
  wire signed [16-1:0] _cond_data_554;
  assign _cond_data_554 = (_eq_data_552)? _cond_data_491 : 1'sd0;
  wire signed [16-1:0] _cond_data_558;
  assign _cond_data_558 = (_eq_data_556)? _cond_data_461 : _cond_data_554;
  wire signed [16-1:0] _cond_data_561;
  assign _cond_data_561 = (_eq_data_559)? _cond_data_431 : _cond_data_558;
  wire signed [16-1:0] _cond_data_564;
  assign _cond_data_564 = (_eq_data_562)? _cond_data_431 : 1'sd0;
  wire signed [16-1:0] _cond_data_568;
  assign _cond_data_568 = (_eq_data_566)? _cond_data_491 : _cond_data_564;
  wire signed [16-1:0] _cond_data_571;
  assign _cond_data_571 = (_eq_data_569)? _cond_data_461 : _cond_data_568;
  wire signed [16-1:0] _cond_data_574;
  assign _cond_data_574 = (_eq_data_572)? _cond_data_461 : 1'sd0;
  wire signed [16-1:0] _cond_data_578;
  assign _cond_data_578 = (_eq_data_576)? _cond_data_431 : _cond_data_574;
  wire signed [16-1:0] _cond_data_581;
  assign _cond_data_581 = (_eq_data_579)? _cond_data_491 : _cond_data_578;
  wire signed [16-1:0] _reinterpretcast_src_618;
  assign _reinterpretcast_src_618 = _cond_data_501;
  wire signed [16-1:0] _reinterpretcast_data_618;
  assign _reinterpretcast_data_618 = _reinterpretcast_src_618;
  wire signed [16-1:0] _reinterpretcast_src_619;
  assign _reinterpretcast_src_619 = _cond_data_531;
  wire signed [16-1:0] _reinterpretcast_data_619;
  assign _reinterpretcast_data_619 = _reinterpretcast_src_619;
  wire signed [16-1:0] _reinterpretcast_src_620;
  assign _reinterpretcast_src_620 = _cond_data_561;
  wire signed [16-1:0] _reinterpretcast_data_620;
  assign _reinterpretcast_data_620 = _reinterpretcast_src_620;
  wire signed [16-1:0] _reinterpretcast_src_621;
  assign _reinterpretcast_src_621 = _cond_data_511;
  wire signed [16-1:0] _reinterpretcast_data_621;
  assign _reinterpretcast_data_621 = _reinterpretcast_src_621;
  wire signed [16-1:0] _reinterpretcast_src_622;
  assign _reinterpretcast_src_622 = _cond_data_541;
  wire signed [16-1:0] _reinterpretcast_data_622;
  assign _reinterpretcast_data_622 = _reinterpretcast_src_622;
  wire signed [16-1:0] _reinterpretcast_src_623;
  assign _reinterpretcast_src_623 = _cond_data_571;
  wire signed [16-1:0] _reinterpretcast_data_623;
  assign _reinterpretcast_data_623 = _reinterpretcast_src_623;
  wire signed [16-1:0] _reinterpretcast_src_624;
  assign _reinterpretcast_src_624 = _cond_data_521;
  wire signed [16-1:0] _reinterpretcast_data_624;
  assign _reinterpretcast_data_624 = _reinterpretcast_src_624;
  wire signed [16-1:0] _reinterpretcast_src_625;
  assign _reinterpretcast_src_625 = _cond_data_551;
  wire signed [16-1:0] _reinterpretcast_data_625;
  assign _reinterpretcast_data_625 = _reinterpretcast_src_625;
  wire signed [16-1:0] _reinterpretcast_src_626;
  assign _reinterpretcast_src_626 = _cond_data_581;
  wire signed [16-1:0] _reinterpretcast_data_626;
  assign _reinterpretcast_data_626 = _reinterpretcast_src_626;
  wire signed [16-1:0] _cond_data_700;
  assign _cond_data_700 = (__delay_data_1263_pointer_681)? 1'sd0 : _reinterpretcast_data_618;
  wire signed [16-1:0] _cond_data_702;
  assign _cond_data_702 = (__delay_data_1265_pointer_683)? 1'sd0 : _reinterpretcast_data_619;
  wire signed [16-1:0] _cond_data_704;
  assign _cond_data_704 = (__delay_data_1267_pointer_685)? 1'sd0 : _reinterpretcast_data_620;
  wire signed [16-1:0] _cond_data_706;
  assign _cond_data_706 = (__delay_data_1269_pointer_687)? 1'sd0 : _reinterpretcast_data_621;
  wire signed [16-1:0] _cond_data_708;
  assign _cond_data_708 = (__delay_data_1271_pointer_689)? 1'sd0 : _reinterpretcast_data_622;
  wire signed [16-1:0] _cond_data_710;
  assign _cond_data_710 = (__delay_data_1273_pointer_691)? 1'sd0 : _reinterpretcast_data_623;
  wire signed [16-1:0] _cond_data_712;
  assign _cond_data_712 = (__delay_data_1275_pointer_693)? 1'sd0 : _reinterpretcast_data_624;
  wire signed [16-1:0] _cond_data_714;
  assign _cond_data_714 = (__delay_data_1277_pointer_695)? 1'sd0 : _reinterpretcast_data_625;
  wire signed [16-1:0] _cond_data_716;
  assign _cond_data_716 = (__delay_data_1279_pointer_697)? 1'sd0 : _reinterpretcast_data_626;
  reg signed [16-1:0] __variable_wdata_136;
  assign mul_8_x_data = __variable_wdata_136;
  reg signed [16-1:0] __variable_wdata_137;
  assign mul_8_y_data = __variable_wdata_137;
  reg [5-1:0] __variable_wdata_138;
  assign mul_8_rshift_data = __variable_wdata_138;
  reg signed [16-1:0] __variable_wdata_157;
  assign mul_9_x_data = __variable_wdata_157;
  reg signed [16-1:0] __variable_wdata_158;
  assign mul_9_y_data = __variable_wdata_158;
  reg [5-1:0] __variable_wdata_159;
  assign mul_9_rshift_data = __variable_wdata_159;
  reg signed [16-1:0] __variable_wdata_178;
  assign mul_10_x_data = __variable_wdata_178;
  reg signed [16-1:0] __variable_wdata_179;
  assign mul_10_y_data = __variable_wdata_179;
  reg [5-1:0] __variable_wdata_180;
  assign mul_10_rshift_data = __variable_wdata_180;
  reg signed [16-1:0] __variable_wdata_199;
  assign mul_11_x_data = __variable_wdata_199;
  reg signed [16-1:0] __variable_wdata_200;
  assign mul_11_y_data = __variable_wdata_200;
  reg [5-1:0] __variable_wdata_201;
  assign mul_11_rshift_data = __variable_wdata_201;
  reg signed [16-1:0] __variable_wdata_220;
  assign mul_12_x_data = __variable_wdata_220;
  reg signed [16-1:0] __variable_wdata_221;
  assign mul_12_y_data = __variable_wdata_221;
  reg [5-1:0] __variable_wdata_222;
  assign mul_12_rshift_data = __variable_wdata_222;
  assign _mul_12_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_12_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_12_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_241;
  assign mul_13_x_data = __variable_wdata_241;
  reg signed [16-1:0] __variable_wdata_242;
  assign mul_13_y_data = __variable_wdata_242;
  reg [5-1:0] __variable_wdata_243;
  assign mul_13_rshift_data = __variable_wdata_243;
  assign _mul_13_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_13_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_13_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_262;
  assign mul_14_x_data = __variable_wdata_262;
  reg signed [16-1:0] __variable_wdata_263;
  assign mul_14_y_data = __variable_wdata_263;
  reg [5-1:0] __variable_wdata_264;
  assign mul_14_rshift_data = __variable_wdata_264;
  assign _mul_14_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_14_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_14_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_283;
  assign mul_15_x_data = __variable_wdata_283;
  reg signed [16-1:0] __variable_wdata_284;
  assign mul_15_y_data = __variable_wdata_284;
  reg [5-1:0] __variable_wdata_285;
  assign mul_15_rshift_data = __variable_wdata_285;
  assign _mul_15_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_15_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_15_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_304;
  assign mul_16_x_data = __variable_wdata_304;
  reg signed [16-1:0] __variable_wdata_305;
  assign mul_16_y_data = __variable_wdata_305;
  reg [5-1:0] __variable_wdata_306;
  assign mul_16_rshift_data = __variable_wdata_306;
  assign _mul_16_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_16_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_16_stream_internal_oready;
  reg [1-1:0] __delay_data_1282__delay_1281__variable_344;
  reg [16-1:0] __delay_data_1294_plus_902;
  reg [8-1:0] __delay_data_1307__delay_1306__variable_339;
  reg signed [16-1:0] __delay_data_1320__delay_1319_cond_360;
  reg signed [16-1:0] __delay_data_1339__delay_1338_cond_367;
  reg [16-1:0] __delay_data_1358_plus_921;
  reg [1-1:0] __delay_data_1283__delay_1282__delay_1281__variable_344;
  reg [16-1:0] __delay_data_1295__delay_1294_plus_902;
  reg [8-1:0] __delay_data_1308__delay_1307__delay_1306__variable_339;
  reg signed [16-1:0] __delay_data_1321__delay_1320__delay_1319_cond_360;
  reg signed [16-1:0] __delay_data_1340__delay_1339__delay_1338_cond_367;
  reg [16-1:0] __delay_data_1359__delay_1358_plus_921;
  reg [1-1:0] __delay_data_1284__delay_1283__delay_1282____variable_344;
  reg [16-1:0] __delay_data_1296__delay_1295__delay_1294_plus_902;
  reg [8-1:0] __delay_data_1309__delay_1308__delay_1307____variable_339;
  reg signed [16-1:0] __delay_data_1322__delay_1321__delay_1320__delay_1319_cond_360;
  reg signed [16-1:0] __delay_data_1341__delay_1340__delay_1339__delay_1338_cond_367;
  reg [16-1:0] __delay_data_1360__delay_1359__delay_1358_plus_921;
  reg [1-1:0] __delay_data_1285__delay_1284__delay_1283____variable_344;
  reg [16-1:0] __delay_data_1297__delay_1296__delay_1295__delay_1294_plus_902;
  reg [8-1:0] __delay_data_1310__delay_1309__delay_1308____variable_339;
  reg signed [16-1:0] __delay_data_1323__delay_1322__delay_1321__delay_1320___cond_360;
  reg signed [16-1:0] __delay_data_1342__delay_1341__delay_1340__delay_1339___cond_367;
  reg [16-1:0] __delay_data_1361__delay_1360__delay_1359__delay_1358_plus_921;
  reg [1-1:0] __delay_data_1286__delay_1285__delay_1284____variable_344;
  reg [16-1:0] __delay_data_1298__delay_1297__delay_1296__delay_1295___plus_902;
  reg [8-1:0] __delay_data_1311__delay_1310__delay_1309____variable_339;
  reg signed [16-1:0] __delay_data_1324__delay_1323__delay_1322__delay_1321___cond_360;
  reg signed [16-1:0] __delay_data_1343__delay_1342__delay_1341__delay_1340___cond_367;
  reg [16-1:0] __delay_data_1362__delay_1361__delay_1360__delay_1359___plus_921;
  reg [1-1:0] __delay_data_1287__delay_1286__delay_1285____variable_344;
  reg [16-1:0] __delay_data_1299__delay_1298__delay_1297__delay_1296___plus_902;
  reg [8-1:0] __delay_data_1312__delay_1311__delay_1310____variable_339;
  reg signed [16-1:0] __delay_data_1325__delay_1324__delay_1323__delay_1322___cond_360;
  reg signed [16-1:0] __delay_data_1344__delay_1343__delay_1342__delay_1341___cond_367;
  reg [16-1:0] __delay_data_1363__delay_1362__delay_1361__delay_1360___plus_921;
  reg [1-1:0] __delay_data_1288__delay_1287__delay_1286____variable_344;
  reg [16-1:0] __delay_data_1300__delay_1299__delay_1298__delay_1297___plus_902;
  reg [8-1:0] __delay_data_1313__delay_1312__delay_1311____variable_339;
  reg signed [16-1:0] __delay_data_1326__delay_1325__delay_1324__delay_1323___cond_360;
  reg signed [16-1:0] __delay_data_1345__delay_1344__delay_1343__delay_1342___cond_367;
  reg [16-1:0] __delay_data_1364__delay_1363__delay_1362__delay_1361___plus_921;
  reg [1-1:0] __delay_data_1289__delay_1288__delay_1287____variable_344;
  reg [16-1:0] __delay_data_1301__delay_1300__delay_1299__delay_1298___plus_902;
  reg [8-1:0] __delay_data_1314__delay_1313__delay_1312____variable_339;
  reg signed [16-1:0] __delay_data_1327__delay_1326__delay_1325__delay_1324___cond_360;
  reg signed [16-1:0] __delay_data_1346__delay_1345__delay_1344__delay_1343___cond_367;
  reg [16-1:0] __delay_data_1365__delay_1364__delay_1363__delay_1362___plus_921;
  reg [1-1:0] __delay_data_1290__delay_1289__delay_1288____variable_344;
  reg [16-1:0] __delay_data_1302__delay_1301__delay_1300__delay_1299___plus_902;
  reg [8-1:0] __delay_data_1315__delay_1314__delay_1313____variable_339;
  reg signed [16-1:0] __delay_data_1328__delay_1327__delay_1326__delay_1325___cond_360;
  reg signed [16-1:0] __delay_data_1347__delay_1346__delay_1345__delay_1344___cond_367;
  reg [16-1:0] __delay_data_1366__delay_1365__delay_1364__delay_1363___plus_921;
  wire signed [32-1:0] __substreamoutput_data_735;
  assign __substreamoutput_data_735 = mul_8_z_data;
  wire signed [32-1:0] __substreamoutput_data_754;
  assign __substreamoutput_data_754 = mul_9_z_data;
  wire signed [32-1:0] __substreamoutput_data_773;
  assign __substreamoutput_data_773 = mul_10_z_data;
  wire signed [32-1:0] __substreamoutput_data_792;
  assign __substreamoutput_data_792 = mul_11_z_data;
  wire signed [32-1:0] __substreamoutput_data_811;
  assign __substreamoutput_data_811 = mul_12_z_data;
  wire signed [32-1:0] __substreamoutput_data_830;
  assign __substreamoutput_data_830 = mul_13_z_data;
  wire signed [32-1:0] __substreamoutput_data_849;
  assign __substreamoutput_data_849 = mul_14_z_data;
  wire signed [32-1:0] __substreamoutput_data_868;
  assign __substreamoutput_data_868 = mul_15_z_data;
  wire signed [32-1:0] __substreamoutput_data_887;
  assign __substreamoutput_data_887 = mul_16_z_data;
  reg signed [64-1:0] __variable_wdata_54;
  assign add_tree_5_var0_data = __variable_wdata_54;
  reg signed [64-1:0] __variable_wdata_55;
  assign add_tree_5_var1_data = __variable_wdata_55;
  reg signed [64-1:0] __variable_wdata_56;
  assign add_tree_5_var2_data = __variable_wdata_56;
  reg signed [64-1:0] __variable_wdata_57;
  assign add_tree_5_var3_data = __variable_wdata_57;
  reg signed [64-1:0] __variable_wdata_58;
  assign add_tree_5_var4_data = __variable_wdata_58;
  reg signed [64-1:0] __variable_wdata_59;
  assign add_tree_5_var5_data = __variable_wdata_59;
  reg signed [64-1:0] __variable_wdata_60;
  assign add_tree_5_var6_data = __variable_wdata_60;
  reg signed [64-1:0] __variable_wdata_61;
  assign add_tree_5_var7_data = __variable_wdata_61;
  reg signed [64-1:0] __variable_wdata_62;
  assign add_tree_5_var8_data = __variable_wdata_62;
  assign _add_tree_5_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _add_tree_5_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _add_tree_5_stream_internal_oready;
  reg [1-1:0] __delay_data_1291__delay_1290__delay_1289____variable_344;
  reg [16-1:0] __delay_data_1303__delay_1302__delay_1301__delay_1300___plus_902;
  reg [8-1:0] __delay_data_1316__delay_1315__delay_1314____variable_339;
  reg signed [16-1:0] __delay_data_1329__delay_1328__delay_1327__delay_1326___cond_360;
  reg signed [16-1:0] __delay_data_1348__delay_1347__delay_1346__delay_1345___cond_367;
  reg [16-1:0] __delay_data_1367__delay_1366__delay_1365__delay_1364___plus_921;
  reg [1-1:0] __delay_data_1292__delay_1291__delay_1290____variable_344;
  reg [16-1:0] __delay_data_1304__delay_1303__delay_1302__delay_1301___plus_902;
  reg [8-1:0] __delay_data_1317__delay_1316__delay_1315____variable_339;
  reg signed [16-1:0] __delay_data_1330__delay_1329__delay_1328__delay_1327___cond_360;
  reg signed [16-1:0] __delay_data_1349__delay_1348__delay_1347__delay_1346___cond_367;
  reg [16-1:0] __delay_data_1368__delay_1367__delay_1366__delay_1365___plus_921;
  reg [1-1:0] __delay_data_1293__delay_1292__delay_1291____variable_344;
  reg [16-1:0] __delay_data_1305__delay_1304__delay_1303__delay_1302___plus_902;
  reg [8-1:0] __delay_data_1318__delay_1317__delay_1316____variable_339;
  reg signed [16-1:0] __delay_data_1331__delay_1330__delay_1329__delay_1328___cond_360;
  reg signed [16-1:0] __delay_data_1350__delay_1349__delay_1348__delay_1347___cond_367;
  reg [16-1:0] __delay_data_1369__delay_1368__delay_1367__delay_1366___plus_921;
  wire signed [64-1:0] __substreamoutput_data_889;
  assign __substreamoutput_data_889 = add_tree_5_sum_data;
  reg [1-1:0] __variable_wdata_15;
  assign acc_0__reduce_reset_data = __variable_wdata_15;
  reg signed [64-1:0] __variable_wdata_0;
  assign acc_0_x_data = __variable_wdata_0;
  reg [7-1:0] __variable_wdata_1;
  assign acc_0_rshift_data = __variable_wdata_1;
  reg [32-1:0] __variable_wdata_2;
  assign acc_0_size_data = __variable_wdata_2;
  reg signed [16-1:0] __delay_data_1332__delay_1331__delay_1330__delay_1329___cond_360;
  reg signed [16-1:0] __delay_data_1351__delay_1350__delay_1349__delay_1348___cond_367;
  reg [16-1:0] __delay_data_1370__delay_1369__delay_1368__delay_1367___plus_921;
  reg signed [16-1:0] __delay_data_1333__delay_1332__delay_1331__delay_1330___cond_360;
  reg signed [16-1:0] __delay_data_1352__delay_1351__delay_1350__delay_1349___cond_367;
  reg [16-1:0] __delay_data_1371__delay_1370__delay_1369__delay_1368___plus_921;
  reg signed [16-1:0] __delay_data_1334__delay_1333__delay_1332__delay_1331___cond_360;
  reg signed [16-1:0] __delay_data_1353__delay_1352__delay_1351__delay_1350___cond_367;
  reg [16-1:0] __delay_data_1372__delay_1371__delay_1370__delay_1369___plus_921;
  reg signed [16-1:0] __delay_data_1335__delay_1334__delay_1333__delay_1332___cond_360;
  reg signed [16-1:0] __delay_data_1354__delay_1353__delay_1352__delay_1351___cond_367;
  reg [16-1:0] __delay_data_1373__delay_1372__delay_1371__delay_1370___plus_921;
  reg signed [16-1:0] __delay_data_1336__delay_1335__delay_1334__delay_1333___cond_360;
  reg signed [16-1:0] __delay_data_1355__delay_1354__delay_1353__delay_1352___cond_367;
  reg [16-1:0] __delay_data_1374__delay_1373__delay_1372__delay_1371___plus_921;
  reg signed [16-1:0] __delay_data_1337__delay_1336__delay_1335__delay_1334___cond_360;
  reg signed [16-1:0] __delay_data_1356__delay_1355__delay_1354__delay_1353___cond_367;
  reg [16-1:0] __delay_data_1375__delay_1374__delay_1373__delay_1372___plus_921;
  wire signed [64-1:0] __substreamoutput_data_903;
  assign __substreamoutput_data_903 = acc_0_sum_data;
  wire [1-1:0] __substreamoutput_data_904;
  assign __substreamoutput_data_904 = acc_0_valid_data;
  reg signed [64-1:0] _plus_data_905;
  reg signed [16-1:0] __delay_data_1357__delay_1356__delay_1355__delay_1354___cond_367;
  reg [16-1:0] __delay_data_1376__delay_1375__delay_1374__delay_1373___plus_921;
  reg [1-1:0] __delay_data_1378__substreamoutput_904;
  reg signed [64-1:0] __variable_wdata_68;
  assign mul_rshift_round_clip_6_x_data = __variable_wdata_68;
  reg signed [16-1:0] __variable_wdata_69;
  assign mul_rshift_round_clip_6_y_data = __variable_wdata_69;
  reg [7-1:0] __variable_wdata_70;
  assign mul_rshift_round_clip_6_rshift_data = __variable_wdata_70;
  assign _stream_conv2d_4_stream_internal_oready = ((_stream_conv2d_4_busy)? _mul_rshift_round_clip_6_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _acc_0_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _add_tree_5_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_16_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_15_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_14_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_13_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_12_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_11_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_10_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_9_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_8_stream_internal_oready : 1) && 1)))))))))));
  reg [1-1:0] __delay_data_1379__delay_1378__substreamoutput_904;
  reg [1-1:0] __delay_data_1380__delay_1379__delay_1378__substreamoutput_904;
  reg [1-1:0] __delay_data_1381__delay_1380__delay_1379____substreamoutput_904;
  reg [1-1:0] __delay_data_1382__delay_1381__delay_1380____substreamoutput_904;
  reg [1-1:0] __delay_data_1383__delay_1382__delay_1381____substreamoutput_904;
  reg [1-1:0] __delay_data_1384__delay_1383__delay_1382____substreamoutput_904;
  reg [1-1:0] __delay_data_1385__delay_1384__delay_1383____substreamoutput_904;
  reg [1-1:0] __delay_data_1386__delay_1385__delay_1384____substreamoutput_904;
  reg [1-1:0] __delay_data_1387__delay_1386__delay_1385____substreamoutput_904;
  wire signed [16-1:0] __substreamoutput_data_922;
  assign __substreamoutput_data_922 = mul_rshift_round_clip_6_z_data;
  reg [1-1:0] _greaterthan_data_924;
  reg signed [16-1:0] __delay_data_1377__substreamoutput_922;
  reg [1-1:0] __delay_data_1388__delay_1387__delay_1386____substreamoutput_904;
  reg signed [16-1:0] _cond_data_926;
  reg [1-1:0] __delay_data_1389__delay_1388__delay_1387____substreamoutput_904;
  wire signed [16-1:0] _reinterpretcast_src_927;
  assign _reinterpretcast_src_927 = _cond_data_926;
  wire signed [16-1:0] _reinterpretcast_data_927;
  assign _reinterpretcast_data_927 = _reinterpretcast_src_927;
  wire signed [16-1:0] stream_conv2d_4_sink_50_data;
  assign stream_conv2d_4_sink_50_data = _reinterpretcast_data_927;
  wire [1-1:0] stream_conv2d_4_sink_51_data;
  assign stream_conv2d_4_sink_51_data = __delay_data_1389__delay_1388__delay_1387____substreamoutput_904;
  wire _set_flag_328;
  assign _set_flag_328 = conv2d_4_comp_fsm == 3;
  reg [8-1:0] __variable_wdata_339;
  assign stream_conv2d_4_parameter_0_data = __variable_wdata_339;
  wire _set_flag_329;
  assign _set_flag_329 = conv2d_4_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_340;
  assign stream_conv2d_4_parameter_1_data = __variable_wdata_340;
  wire _set_flag_330;
  assign _set_flag_330 = conv2d_4_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_341;
  assign stream_conv2d_4_parameter_2_data = __variable_wdata_341;
  wire _set_flag_331;
  assign _set_flag_331 = conv2d_4_comp_fsm == 3;
  reg [9-1:0] __variable_wdata_342;
  assign stream_conv2d_4_parameter_3_data = __variable_wdata_342;
  wire _set_flag_332;
  assign _set_flag_332 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_343;
  assign stream_conv2d_4_parameter_4_data = __variable_wdata_343;
  wire _set_flag_333;
  assign _set_flag_333 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_354;
  assign stream_conv2d_4_parameter_6_data = __variable_wdata_354;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_buf_3;
  wire _set_flag_334;
  assign _set_flag_334 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_335;
  assign read_rtl_bank_335 = _stream_conv2d_4_source_7_source_ram_raddr;
  reg [1-1:0] _tmp_336;
  assign ram_w16_l512_id1_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1))? _stream_conv2d_4_source_7_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id1_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_337 = 1;
  wire [_tmp_337-1:0] _tmp_338;
  assign _tmp_338 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1);
  reg [_tmp_337-1:0] __tmp_338_1;
  assign ram_w16_l512_id1_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1))? _stream_conv2d_4_source_7_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id1_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_339 = 1;
  wire [_tmp_339-1:0] _tmp_340;
  assign _tmp_340 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1);
  reg [_tmp_339-1:0] __tmp_340_1;
  wire signed [16-1:0] read_rtl_rdata_341;
  wire read_rtl_rvalid_342;
  assign read_rtl_rdata_341 = (_tmp_336 == 0)? ram_w16_l512_id1_0_0_rdata : 
                              (_tmp_336 == 1)? ram_w16_l512_id1_1_0_rdata : 0;
  assign read_rtl_rvalid_342 = __tmp_338_1;
  assign _stream_conv2d_4_source_7_source_ram_rdata = (_stream_conv2d_4_source_7_source_sel == 1)? read_rtl_rdata_341 : 'hx;
  reg [16-1:0] __variable_wdata_355;
  assign stream_conv2d_4_source_7_data = __variable_wdata_355;
  reg [32-1:0] _stream_conv2d_4_source_7_source_pat_fsm_0;
  localparam _stream_conv2d_4_source_7_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_7_source_pat_all_offset;
  assign _stream_conv2d_4_source_7_source_pat_all_offset = _stream_conv2d_4_source_7_source_offset_buf + _source_stream_conv2d_4_source_7_pat_cur_offset_0 + _source_stream_conv2d_4_source_7_pat_cur_offset_1 + _source_stream_conv2d_4_source_7_pat_cur_offset_2 + _source_stream_conv2d_4_source_7_pat_cur_offset_3;
  wire _set_flag_343;
  assign _set_flag_343 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_361;
  assign stream_conv2d_4_parameter_8_data = __variable_wdata_361;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_buf_3;
  wire _set_flag_344;
  assign _set_flag_344 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_345;
  assign read_rtl_bank_345 = _stream_conv2d_4_source_9_source_ram_raddr;
  reg [1-1:0] _tmp_346;
  assign ram_w16_l512_id2_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2))? _stream_conv2d_4_source_9_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id2_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_347 = 1;
  wire [_tmp_347-1:0] _tmp_348;
  assign _tmp_348 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2);
  reg [_tmp_347-1:0] __tmp_348_1;
  assign ram_w16_l512_id2_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2))? _stream_conv2d_4_source_9_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id2_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_349 = 1;
  wire [_tmp_349-1:0] _tmp_350;
  assign _tmp_350 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2);
  reg [_tmp_349-1:0] __tmp_350_1;
  wire signed [16-1:0] read_rtl_rdata_351;
  wire read_rtl_rvalid_352;
  assign read_rtl_rdata_351 = (_tmp_346 == 0)? ram_w16_l512_id2_0_0_rdata : 
                              (_tmp_346 == 1)? ram_w16_l512_id2_1_0_rdata : 0;
  assign read_rtl_rvalid_352 = __tmp_348_1;
  assign _stream_conv2d_4_source_9_source_ram_rdata = (_stream_conv2d_4_source_9_source_sel == 2)? read_rtl_rdata_351 : 'hx;
  reg [16-1:0] __variable_wdata_362;
  assign stream_conv2d_4_source_9_data = __variable_wdata_362;
  reg [32-1:0] _stream_conv2d_4_source_9_source_pat_fsm_1;
  localparam _stream_conv2d_4_source_9_source_pat_fsm_1_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_9_source_pat_all_offset;
  assign _stream_conv2d_4_source_9_source_pat_all_offset = _stream_conv2d_4_source_9_source_offset_buf + _source_stream_conv2d_4_source_9_pat_cur_offset_0 + _source_stream_conv2d_4_source_9_pat_cur_offset_1 + _source_stream_conv2d_4_source_9_pat_cur_offset_2 + _source_stream_conv2d_4_source_9_pat_cur_offset_3;
  wire _set_flag_353;
  assign _set_flag_353 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_368;
  assign stream_conv2d_4_parameter_10_data = __variable_wdata_368;
  wire _set_flag_354;
  assign _set_flag_354 = conv2d_4_comp_fsm == 3;
  reg [16-1:0] __variable_wdata_369;
  assign stream_conv2d_4_source_11_data = __variable_wdata_369;
  wire _set_flag_355;
  assign _set_flag_355 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_375;
  assign stream_conv2d_4_parameter_12_data = __variable_wdata_375;
  wire _set_flag_356;
  assign _set_flag_356 = conv2d_4_comp_fsm == 3;
  reg [16-1:0] __variable_wdata_376;
  assign stream_conv2d_4_source_13_data = __variable_wdata_376;
  wire _set_flag_357;
  assign _set_flag_357 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_382;
  assign stream_conv2d_4_parameter_14_data = __variable_wdata_382;
  wire _set_flag_358;
  assign _set_flag_358 = conv2d_4_comp_fsm == 3;
  reg [16-1:0] __variable_wdata_383;
  assign stream_conv2d_4_source_15_data = __variable_wdata_383;
  wire _set_flag_359;
  assign _set_flag_359 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_389;
  assign stream_conv2d_4_parameter_16_data = __variable_wdata_389;
  wire _set_flag_360;
  assign _set_flag_360 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_390;
  assign stream_conv2d_4_parameter_17_data = __variable_wdata_390;
  wire _set_flag_361;
  assign _set_flag_361 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_391;
  assign stream_conv2d_4_parameter_18_data = __variable_wdata_391;
  wire _set_flag_362;
  assign _set_flag_362 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_392;
  assign stream_conv2d_4_parameter_19_data = __variable_wdata_392;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_buf_3;
  wire _set_flag_363;
  assign _set_flag_363 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_364;
  assign read_rtl_bank_364 = _stream_conv2d_4_source_20_source_ram_raddr;
  reg [1-1:0] _tmp_365;
  localparam _tmp_366 = 1;
  wire [_tmp_366-1:0] _tmp_367;
  assign _tmp_367 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3);
  reg [_tmp_366-1:0] __tmp_367_1;
  localparam _tmp_368 = 1;
  wire [_tmp_368-1:0] _tmp_369;
  assign _tmp_369 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3);
  reg [_tmp_368-1:0] __tmp_369_1;
  wire signed [16-1:0] read_rtl_rdata_370;
  wire read_rtl_rvalid_371;
  assign read_rtl_rdata_370 = (_tmp_365 == 0)? ram_w16_l1024_id0_0_0_rdata : 
                              (_tmp_365 == 1)? ram_w16_l1024_id0_1_0_rdata : 0;
  assign read_rtl_rvalid_371 = __tmp_367_1;
  assign _stream_conv2d_4_source_20_source_ram_rdata = (_stream_conv2d_4_source_20_source_sel == 3)? read_rtl_rdata_370 : 'hx;
  reg [16-1:0] __variable_wdata_393;
  assign stream_conv2d_4_source_20_data = __variable_wdata_393;
  reg [32-1:0] _stream_conv2d_4_source_20_source_pat_fsm_2;
  localparam _stream_conv2d_4_source_20_source_pat_fsm_2_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_20_source_pat_all_offset;
  assign _stream_conv2d_4_source_20_source_pat_all_offset = _stream_conv2d_4_source_20_source_offset_buf + _source_stream_conv2d_4_source_20_pat_cur_offset_0 + _source_stream_conv2d_4_source_20_pat_cur_offset_1 + _source_stream_conv2d_4_source_20_pat_cur_offset_2 + _source_stream_conv2d_4_source_20_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_buf_3;
  wire _set_flag_372;
  assign _set_flag_372 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_373;
  assign read_rtl_bank_373 = _stream_conv2d_4_source_21_source_ram_raddr;
  reg [1-1:0] _tmp_374;
  localparam _tmp_375 = 1;
  wire [_tmp_375-1:0] _tmp_376;
  assign _tmp_376 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4);
  reg [_tmp_375-1:0] __tmp_376_1;
  localparam _tmp_377 = 1;
  wire [_tmp_377-1:0] _tmp_378;
  assign _tmp_378 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4);
  reg [_tmp_377-1:0] __tmp_378_1;
  wire signed [16-1:0] read_rtl_rdata_379;
  wire read_rtl_rvalid_380;
  assign read_rtl_rdata_379 = (_tmp_374 == 0)? ram_w16_l1024_id1_0_0_rdata : 
                              (_tmp_374 == 1)? ram_w16_l1024_id1_1_0_rdata : 0;
  assign read_rtl_rvalid_380 = __tmp_376_1;
  assign _stream_conv2d_4_source_21_source_ram_rdata = (_stream_conv2d_4_source_21_source_sel == 4)? read_rtl_rdata_379 : 'hx;
  reg [16-1:0] __variable_wdata_394;
  assign stream_conv2d_4_source_21_data = __variable_wdata_394;
  reg [32-1:0] _stream_conv2d_4_source_21_source_pat_fsm_3;
  localparam _stream_conv2d_4_source_21_source_pat_fsm_3_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_21_source_pat_all_offset;
  assign _stream_conv2d_4_source_21_source_pat_all_offset = _stream_conv2d_4_source_21_source_offset_buf + _source_stream_conv2d_4_source_21_pat_cur_offset_0 + _source_stream_conv2d_4_source_21_pat_cur_offset_1 + _source_stream_conv2d_4_source_21_pat_cur_offset_2 + _source_stream_conv2d_4_source_21_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_buf_3;
  wire _set_flag_381;
  assign _set_flag_381 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_382;
  assign read_rtl_bank_382 = _stream_conv2d_4_source_22_source_ram_raddr;
  reg [1-1:0] _tmp_383;
  assign ram_w16_l1024_id2_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5))? _stream_conv2d_4_source_22_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id2_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5))? 1'd1 : 0;
  localparam _tmp_384 = 1;
  wire [_tmp_384-1:0] _tmp_385;
  assign _tmp_385 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5);
  reg [_tmp_384-1:0] __tmp_385_1;
  assign ram_w16_l1024_id2_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5))? _stream_conv2d_4_source_22_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id2_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5))? 1'd1 : 0;
  localparam _tmp_386 = 1;
  wire [_tmp_386-1:0] _tmp_387;
  assign _tmp_387 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5);
  reg [_tmp_386-1:0] __tmp_387_1;
  wire signed [16-1:0] read_rtl_rdata_388;
  wire read_rtl_rvalid_389;
  assign read_rtl_rdata_388 = (_tmp_383 == 0)? ram_w16_l1024_id2_0_0_rdata : 
                              (_tmp_383 == 1)? ram_w16_l1024_id2_1_0_rdata : 0;
  assign read_rtl_rvalid_389 = __tmp_385_1;
  assign _stream_conv2d_4_source_22_source_ram_rdata = (_stream_conv2d_4_source_22_source_sel == 5)? read_rtl_rdata_388 : 'hx;
  reg [16-1:0] __variable_wdata_395;
  assign stream_conv2d_4_source_22_data = __variable_wdata_395;
  reg [32-1:0] _stream_conv2d_4_source_22_source_pat_fsm_4;
  localparam _stream_conv2d_4_source_22_source_pat_fsm_4_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_22_source_pat_all_offset;
  assign _stream_conv2d_4_source_22_source_pat_all_offset = _stream_conv2d_4_source_22_source_offset_buf + _source_stream_conv2d_4_source_22_pat_cur_offset_0 + _source_stream_conv2d_4_source_22_pat_cur_offset_1 + _source_stream_conv2d_4_source_22_pat_cur_offset_2 + _source_stream_conv2d_4_source_22_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_buf_3;
  wire _set_flag_390;
  assign _set_flag_390 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_391;
  assign read_rtl_bank_391 = _stream_conv2d_4_source_23_source_ram_raddr;
  reg [1-1:0] _tmp_392;
  assign ram_w16_l1024_id3_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6))? _stream_conv2d_4_source_23_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id3_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6))? 1'd1 : 0;
  localparam _tmp_393 = 1;
  wire [_tmp_393-1:0] _tmp_394;
  assign _tmp_394 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6);
  reg [_tmp_393-1:0] __tmp_394_1;
  assign ram_w16_l1024_id3_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6))? _stream_conv2d_4_source_23_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id3_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6))? 1'd1 : 0;
  localparam _tmp_395 = 1;
  wire [_tmp_395-1:0] _tmp_396;
  assign _tmp_396 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6);
  reg [_tmp_395-1:0] __tmp_396_1;
  wire signed [16-1:0] read_rtl_rdata_397;
  wire read_rtl_rvalid_398;
  assign read_rtl_rdata_397 = (_tmp_392 == 0)? ram_w16_l1024_id3_0_0_rdata : 
                              (_tmp_392 == 1)? ram_w16_l1024_id3_1_0_rdata : 0;
  assign read_rtl_rvalid_398 = __tmp_394_1;
  assign _stream_conv2d_4_source_23_source_ram_rdata = (_stream_conv2d_4_source_23_source_sel == 6)? read_rtl_rdata_397 : 'hx;
  reg [16-1:0] __variable_wdata_396;
  assign stream_conv2d_4_source_23_data = __variable_wdata_396;
  reg [32-1:0] _stream_conv2d_4_source_23_source_pat_fsm_5;
  localparam _stream_conv2d_4_source_23_source_pat_fsm_5_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_23_source_pat_all_offset;
  assign _stream_conv2d_4_source_23_source_pat_all_offset = _stream_conv2d_4_source_23_source_offset_buf + _source_stream_conv2d_4_source_23_pat_cur_offset_0 + _source_stream_conv2d_4_source_23_pat_cur_offset_1 + _source_stream_conv2d_4_source_23_pat_cur_offset_2 + _source_stream_conv2d_4_source_23_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_buf_3;
  wire _set_flag_399;
  assign _set_flag_399 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_400;
  assign read_rtl_bank_400 = _stream_conv2d_4_source_24_source_ram_raddr;
  reg [1-1:0] _tmp_401;
  assign ram_w16_l1024_id4_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7))? _stream_conv2d_4_source_24_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id4_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7))? 1'd1 : 0;
  localparam _tmp_402 = 1;
  wire [_tmp_402-1:0] _tmp_403;
  assign _tmp_403 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7);
  reg [_tmp_402-1:0] __tmp_403_1;
  assign ram_w16_l1024_id4_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7))? _stream_conv2d_4_source_24_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id4_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7))? 1'd1 : 0;
  localparam _tmp_404 = 1;
  wire [_tmp_404-1:0] _tmp_405;
  assign _tmp_405 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7);
  reg [_tmp_404-1:0] __tmp_405_1;
  wire signed [16-1:0] read_rtl_rdata_406;
  wire read_rtl_rvalid_407;
  assign read_rtl_rdata_406 = (_tmp_401 == 0)? ram_w16_l1024_id4_0_0_rdata : 
                              (_tmp_401 == 1)? ram_w16_l1024_id4_1_0_rdata : 0;
  assign read_rtl_rvalid_407 = __tmp_403_1;
  assign _stream_conv2d_4_source_24_source_ram_rdata = (_stream_conv2d_4_source_24_source_sel == 7)? read_rtl_rdata_406 : 'hx;
  reg [16-1:0] __variable_wdata_397;
  assign stream_conv2d_4_source_24_data = __variable_wdata_397;
  reg [32-1:0] _stream_conv2d_4_source_24_source_pat_fsm_6;
  localparam _stream_conv2d_4_source_24_source_pat_fsm_6_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_24_source_pat_all_offset;
  assign _stream_conv2d_4_source_24_source_pat_all_offset = _stream_conv2d_4_source_24_source_offset_buf + _source_stream_conv2d_4_source_24_pat_cur_offset_0 + _source_stream_conv2d_4_source_24_pat_cur_offset_1 + _source_stream_conv2d_4_source_24_pat_cur_offset_2 + _source_stream_conv2d_4_source_24_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_buf_3;
  wire _set_flag_408;
  assign _set_flag_408 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_409;
  assign read_rtl_bank_409 = _stream_conv2d_4_source_25_source_ram_raddr;
  reg [1-1:0] _tmp_410;
  assign ram_w16_l1024_id5_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8))? _stream_conv2d_4_source_25_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id5_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8))? 1'd1 : 0;
  localparam _tmp_411 = 1;
  wire [_tmp_411-1:0] _tmp_412;
  assign _tmp_412 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8);
  reg [_tmp_411-1:0] __tmp_412_1;
  assign ram_w16_l1024_id5_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8))? _stream_conv2d_4_source_25_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id5_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8))? 1'd1 : 0;
  localparam _tmp_413 = 1;
  wire [_tmp_413-1:0] _tmp_414;
  assign _tmp_414 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8);
  reg [_tmp_413-1:0] __tmp_414_1;
  wire signed [16-1:0] read_rtl_rdata_415;
  wire read_rtl_rvalid_416;
  assign read_rtl_rdata_415 = (_tmp_410 == 0)? ram_w16_l1024_id5_0_0_rdata : 
                              (_tmp_410 == 1)? ram_w16_l1024_id5_1_0_rdata : 0;
  assign read_rtl_rvalid_416 = __tmp_412_1;
  assign _stream_conv2d_4_source_25_source_ram_rdata = (_stream_conv2d_4_source_25_source_sel == 8)? read_rtl_rdata_415 : 'hx;
  reg [16-1:0] __variable_wdata_398;
  assign stream_conv2d_4_source_25_data = __variable_wdata_398;
  reg [32-1:0] _stream_conv2d_4_source_25_source_pat_fsm_7;
  localparam _stream_conv2d_4_source_25_source_pat_fsm_7_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_25_source_pat_all_offset;
  assign _stream_conv2d_4_source_25_source_pat_all_offset = _stream_conv2d_4_source_25_source_offset_buf + _source_stream_conv2d_4_source_25_pat_cur_offset_0 + _source_stream_conv2d_4_source_25_pat_cur_offset_1 + _source_stream_conv2d_4_source_25_pat_cur_offset_2 + _source_stream_conv2d_4_source_25_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_buf_3;
  wire _set_flag_417;
  assign _set_flag_417 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_418;
  assign read_rtl_bank_418 = _stream_conv2d_4_source_26_source_ram_raddr;
  reg [1-1:0] _tmp_419;
  assign ram_w16_l1024_id6_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9))? _stream_conv2d_4_source_26_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id6_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9))? 1'd1 : 0;
  localparam _tmp_420 = 1;
  wire [_tmp_420-1:0] _tmp_421;
  assign _tmp_421 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9);
  reg [_tmp_420-1:0] __tmp_421_1;
  assign ram_w16_l1024_id6_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9))? _stream_conv2d_4_source_26_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id6_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9))? 1'd1 : 0;
  localparam _tmp_422 = 1;
  wire [_tmp_422-1:0] _tmp_423;
  assign _tmp_423 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9);
  reg [_tmp_422-1:0] __tmp_423_1;
  wire signed [16-1:0] read_rtl_rdata_424;
  wire read_rtl_rvalid_425;
  assign read_rtl_rdata_424 = (_tmp_419 == 0)? ram_w16_l1024_id6_0_0_rdata : 
                              (_tmp_419 == 1)? ram_w16_l1024_id6_1_0_rdata : 0;
  assign read_rtl_rvalid_425 = __tmp_421_1;
  assign _stream_conv2d_4_source_26_source_ram_rdata = (_stream_conv2d_4_source_26_source_sel == 9)? read_rtl_rdata_424 : 'hx;
  reg [16-1:0] __variable_wdata_399;
  assign stream_conv2d_4_source_26_data = __variable_wdata_399;
  reg [32-1:0] _stream_conv2d_4_source_26_source_pat_fsm_8;
  localparam _stream_conv2d_4_source_26_source_pat_fsm_8_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_26_source_pat_all_offset;
  assign _stream_conv2d_4_source_26_source_pat_all_offset = _stream_conv2d_4_source_26_source_offset_buf + _source_stream_conv2d_4_source_26_pat_cur_offset_0 + _source_stream_conv2d_4_source_26_pat_cur_offset_1 + _source_stream_conv2d_4_source_26_pat_cur_offset_2 + _source_stream_conv2d_4_source_26_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_buf_3;
  wire _set_flag_426;
  assign _set_flag_426 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_427;
  assign read_rtl_bank_427 = _stream_conv2d_4_source_27_source_ram_raddr;
  reg [1-1:0] _tmp_428;
  assign ram_w16_l1024_id7_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10))? _stream_conv2d_4_source_27_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id7_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10))? 1'd1 : 0;
  localparam _tmp_429 = 1;
  wire [_tmp_429-1:0] _tmp_430;
  assign _tmp_430 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10);
  reg [_tmp_429-1:0] __tmp_430_1;
  assign ram_w16_l1024_id7_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10))? _stream_conv2d_4_source_27_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id7_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10))? 1'd1 : 0;
  localparam _tmp_431 = 1;
  wire [_tmp_431-1:0] _tmp_432;
  assign _tmp_432 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10);
  reg [_tmp_431-1:0] __tmp_432_1;
  wire signed [16-1:0] read_rtl_rdata_433;
  wire read_rtl_rvalid_434;
  assign read_rtl_rdata_433 = (_tmp_428 == 0)? ram_w16_l1024_id7_0_0_rdata : 
                              (_tmp_428 == 1)? ram_w16_l1024_id7_1_0_rdata : 0;
  assign read_rtl_rvalid_434 = __tmp_430_1;
  assign _stream_conv2d_4_source_27_source_ram_rdata = (_stream_conv2d_4_source_27_source_sel == 10)? read_rtl_rdata_433 : 'hx;
  reg [16-1:0] __variable_wdata_400;
  assign stream_conv2d_4_source_27_data = __variable_wdata_400;
  reg [32-1:0] _stream_conv2d_4_source_27_source_pat_fsm_9;
  localparam _stream_conv2d_4_source_27_source_pat_fsm_9_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_27_source_pat_all_offset;
  assign _stream_conv2d_4_source_27_source_pat_all_offset = _stream_conv2d_4_source_27_source_offset_buf + _source_stream_conv2d_4_source_27_pat_cur_offset_0 + _source_stream_conv2d_4_source_27_pat_cur_offset_1 + _source_stream_conv2d_4_source_27_pat_cur_offset_2 + _source_stream_conv2d_4_source_27_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_buf_3;
  wire _set_flag_435;
  assign _set_flag_435 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_436;
  assign read_rtl_bank_436 = _stream_conv2d_4_source_28_source_ram_raddr;
  reg [1-1:0] _tmp_437;
  assign ram_w16_l1024_id8_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11))? _stream_conv2d_4_source_28_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id8_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11))? 1'd1 : 0;
  localparam _tmp_438 = 1;
  wire [_tmp_438-1:0] _tmp_439;
  assign _tmp_439 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11);
  reg [_tmp_438-1:0] __tmp_439_1;
  assign ram_w16_l1024_id8_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11))? _stream_conv2d_4_source_28_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id8_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11))? 1'd1 : 0;
  localparam _tmp_440 = 1;
  wire [_tmp_440-1:0] _tmp_441;
  assign _tmp_441 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11);
  reg [_tmp_440-1:0] __tmp_441_1;
  wire signed [16-1:0] read_rtl_rdata_442;
  wire read_rtl_rvalid_443;
  assign read_rtl_rdata_442 = (_tmp_437 == 0)? ram_w16_l1024_id8_0_0_rdata : 
                              (_tmp_437 == 1)? ram_w16_l1024_id8_1_0_rdata : 0;
  assign read_rtl_rvalid_443 = __tmp_439_1;
  assign _stream_conv2d_4_source_28_source_ram_rdata = (_stream_conv2d_4_source_28_source_sel == 11)? read_rtl_rdata_442 : 'hx;
  reg [16-1:0] __variable_wdata_401;
  assign stream_conv2d_4_source_28_data = __variable_wdata_401;
  reg [32-1:0] _stream_conv2d_4_source_28_source_pat_fsm_10;
  localparam _stream_conv2d_4_source_28_source_pat_fsm_10_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_28_source_pat_all_offset;
  assign _stream_conv2d_4_source_28_source_pat_all_offset = _stream_conv2d_4_source_28_source_offset_buf + _source_stream_conv2d_4_source_28_pat_cur_offset_0 + _source_stream_conv2d_4_source_28_pat_cur_offset_1 + _source_stream_conv2d_4_source_28_pat_cur_offset_2 + _source_stream_conv2d_4_source_28_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_buf_3;
  wire _set_flag_444;
  assign _set_flag_444 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_445;
  assign read_rtl_bank_445 = _stream_conv2d_4_source_29_source_ram_raddr;
  reg [1-1:0] _tmp_446;
  assign ram_w16_l512_id3_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12))? _stream_conv2d_4_source_29_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id3_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12))? 1'd1 : 0;
  localparam _tmp_447 = 1;
  wire [_tmp_447-1:0] _tmp_448;
  assign _tmp_448 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12);
  reg [_tmp_447-1:0] __tmp_448_1;
  assign ram_w16_l512_id3_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12))? _stream_conv2d_4_source_29_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id3_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12))? 1'd1 : 0;
  localparam _tmp_449 = 1;
  wire [_tmp_449-1:0] _tmp_450;
  assign _tmp_450 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12);
  reg [_tmp_449-1:0] __tmp_450_1;
  wire signed [16-1:0] read_rtl_rdata_451;
  wire read_rtl_rvalid_452;
  assign read_rtl_rdata_451 = (_tmp_446 == 0)? ram_w16_l512_id3_0_0_rdata : 
                              (_tmp_446 == 1)? ram_w16_l512_id3_1_0_rdata : 0;
  assign read_rtl_rvalid_452 = __tmp_448_1;
  assign _stream_conv2d_4_source_29_source_ram_rdata = (_stream_conv2d_4_source_29_source_sel == 12)? read_rtl_rdata_451 : 'hx;
  reg [16-1:0] __variable_wdata_627;
  assign stream_conv2d_4_source_29_data = __variable_wdata_627;
  reg [32-1:0] _stream_conv2d_4_source_29_source_pat_fsm_11;
  localparam _stream_conv2d_4_source_29_source_pat_fsm_11_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_29_source_pat_all_offset;
  assign _stream_conv2d_4_source_29_source_pat_all_offset = _stream_conv2d_4_source_29_source_offset_buf + _source_stream_conv2d_4_source_29_pat_cur_offset_0 + _source_stream_conv2d_4_source_29_pat_cur_offset_1 + _source_stream_conv2d_4_source_29_pat_cur_offset_2 + _source_stream_conv2d_4_source_29_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_buf_3;
  wire _set_flag_453;
  assign _set_flag_453 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_454;
  assign read_rtl_bank_454 = _stream_conv2d_4_source_30_source_ram_raddr;
  reg [1-1:0] _tmp_455;
  assign ram_w16_l512_id4_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13))? _stream_conv2d_4_source_30_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id4_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13))? 1'd1 : 0;
  localparam _tmp_456 = 1;
  wire [_tmp_456-1:0] _tmp_457;
  assign _tmp_457 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13);
  reg [_tmp_456-1:0] __tmp_457_1;
  assign ram_w16_l512_id4_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13))? _stream_conv2d_4_source_30_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id4_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13))? 1'd1 : 0;
  localparam _tmp_458 = 1;
  wire [_tmp_458-1:0] _tmp_459;
  assign _tmp_459 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13);
  reg [_tmp_458-1:0] __tmp_459_1;
  wire signed [16-1:0] read_rtl_rdata_460;
  wire read_rtl_rvalid_461;
  assign read_rtl_rdata_460 = (_tmp_455 == 0)? ram_w16_l512_id4_0_0_rdata : 
                              (_tmp_455 == 1)? ram_w16_l512_id4_1_0_rdata : 0;
  assign read_rtl_rvalid_461 = __tmp_457_1;
  assign _stream_conv2d_4_source_30_source_ram_rdata = (_stream_conv2d_4_source_30_source_sel == 13)? read_rtl_rdata_460 : 'hx;
  reg [16-1:0] __variable_wdata_628;
  assign stream_conv2d_4_source_30_data = __variable_wdata_628;
  reg [32-1:0] _stream_conv2d_4_source_30_source_pat_fsm_12;
  localparam _stream_conv2d_4_source_30_source_pat_fsm_12_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_30_source_pat_all_offset;
  assign _stream_conv2d_4_source_30_source_pat_all_offset = _stream_conv2d_4_source_30_source_offset_buf + _source_stream_conv2d_4_source_30_pat_cur_offset_0 + _source_stream_conv2d_4_source_30_pat_cur_offset_1 + _source_stream_conv2d_4_source_30_pat_cur_offset_2 + _source_stream_conv2d_4_source_30_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_buf_3;
  wire _set_flag_462;
  assign _set_flag_462 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_463;
  assign read_rtl_bank_463 = _stream_conv2d_4_source_31_source_ram_raddr;
  reg [1-1:0] _tmp_464;
  assign ram_w16_l512_id5_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14))? _stream_conv2d_4_source_31_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id5_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14))? 1'd1 : 0;
  localparam _tmp_465 = 1;
  wire [_tmp_465-1:0] _tmp_466;
  assign _tmp_466 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14);
  reg [_tmp_465-1:0] __tmp_466_1;
  assign ram_w16_l512_id5_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14))? _stream_conv2d_4_source_31_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id5_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14))? 1'd1 : 0;
  localparam _tmp_467 = 1;
  wire [_tmp_467-1:0] _tmp_468;
  assign _tmp_468 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14);
  reg [_tmp_467-1:0] __tmp_468_1;
  wire signed [16-1:0] read_rtl_rdata_469;
  wire read_rtl_rvalid_470;
  assign read_rtl_rdata_469 = (_tmp_464 == 0)? ram_w16_l512_id5_0_0_rdata : 
                              (_tmp_464 == 1)? ram_w16_l512_id5_1_0_rdata : 0;
  assign read_rtl_rvalid_470 = __tmp_466_1;
  assign _stream_conv2d_4_source_31_source_ram_rdata = (_stream_conv2d_4_source_31_source_sel == 14)? read_rtl_rdata_469 : 'hx;
  reg [16-1:0] __variable_wdata_629;
  assign stream_conv2d_4_source_31_data = __variable_wdata_629;
  reg [32-1:0] _stream_conv2d_4_source_31_source_pat_fsm_13;
  localparam _stream_conv2d_4_source_31_source_pat_fsm_13_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_31_source_pat_all_offset;
  assign _stream_conv2d_4_source_31_source_pat_all_offset = _stream_conv2d_4_source_31_source_offset_buf + _source_stream_conv2d_4_source_31_pat_cur_offset_0 + _source_stream_conv2d_4_source_31_pat_cur_offset_1 + _source_stream_conv2d_4_source_31_pat_cur_offset_2 + _source_stream_conv2d_4_source_31_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_buf_3;
  wire _set_flag_471;
  assign _set_flag_471 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_472;
  assign read_rtl_bank_472 = _stream_conv2d_4_source_32_source_ram_raddr;
  reg [1-1:0] _tmp_473;
  assign ram_w16_l512_id6_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15))? _stream_conv2d_4_source_32_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id6_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15))? 1'd1 : 0;
  localparam _tmp_474 = 1;
  wire [_tmp_474-1:0] _tmp_475;
  assign _tmp_475 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15);
  reg [_tmp_474-1:0] __tmp_475_1;
  assign ram_w16_l512_id6_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15))? _stream_conv2d_4_source_32_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id6_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15))? 1'd1 : 0;
  localparam _tmp_476 = 1;
  wire [_tmp_476-1:0] _tmp_477;
  assign _tmp_477 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15);
  reg [_tmp_476-1:0] __tmp_477_1;
  wire signed [16-1:0] read_rtl_rdata_478;
  wire read_rtl_rvalid_479;
  assign read_rtl_rdata_478 = (_tmp_473 == 0)? ram_w16_l512_id6_0_0_rdata : 
                              (_tmp_473 == 1)? ram_w16_l512_id6_1_0_rdata : 0;
  assign read_rtl_rvalid_479 = __tmp_475_1;
  assign _stream_conv2d_4_source_32_source_ram_rdata = (_stream_conv2d_4_source_32_source_sel == 15)? read_rtl_rdata_478 : 'hx;
  reg [16-1:0] __variable_wdata_630;
  assign stream_conv2d_4_source_32_data = __variable_wdata_630;
  reg [32-1:0] _stream_conv2d_4_source_32_source_pat_fsm_14;
  localparam _stream_conv2d_4_source_32_source_pat_fsm_14_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_32_source_pat_all_offset;
  assign _stream_conv2d_4_source_32_source_pat_all_offset = _stream_conv2d_4_source_32_source_offset_buf + _source_stream_conv2d_4_source_32_pat_cur_offset_0 + _source_stream_conv2d_4_source_32_pat_cur_offset_1 + _source_stream_conv2d_4_source_32_pat_cur_offset_2 + _source_stream_conv2d_4_source_32_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_buf_3;
  wire _set_flag_480;
  assign _set_flag_480 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_481;
  assign read_rtl_bank_481 = _stream_conv2d_4_source_33_source_ram_raddr;
  reg [1-1:0] _tmp_482;
  assign ram_w16_l512_id7_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16))? _stream_conv2d_4_source_33_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id7_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16))? 1'd1 : 0;
  localparam _tmp_483 = 1;
  wire [_tmp_483-1:0] _tmp_484;
  assign _tmp_484 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16);
  reg [_tmp_483-1:0] __tmp_484_1;
  assign ram_w16_l512_id7_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16))? _stream_conv2d_4_source_33_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id7_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16))? 1'd1 : 0;
  localparam _tmp_485 = 1;
  wire [_tmp_485-1:0] _tmp_486;
  assign _tmp_486 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16);
  reg [_tmp_485-1:0] __tmp_486_1;
  wire signed [16-1:0] read_rtl_rdata_487;
  wire read_rtl_rvalid_488;
  assign read_rtl_rdata_487 = (_tmp_482 == 0)? ram_w16_l512_id7_0_0_rdata : 
                              (_tmp_482 == 1)? ram_w16_l512_id7_1_0_rdata : 0;
  assign read_rtl_rvalid_488 = __tmp_484_1;
  assign _stream_conv2d_4_source_33_source_ram_rdata = (_stream_conv2d_4_source_33_source_sel == 16)? read_rtl_rdata_487 : 'hx;
  reg [16-1:0] __variable_wdata_631;
  assign stream_conv2d_4_source_33_data = __variable_wdata_631;
  reg [32-1:0] _stream_conv2d_4_source_33_source_pat_fsm_15;
  localparam _stream_conv2d_4_source_33_source_pat_fsm_15_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_33_source_pat_all_offset;
  assign _stream_conv2d_4_source_33_source_pat_all_offset = _stream_conv2d_4_source_33_source_offset_buf + _source_stream_conv2d_4_source_33_pat_cur_offset_0 + _source_stream_conv2d_4_source_33_pat_cur_offset_1 + _source_stream_conv2d_4_source_33_pat_cur_offset_2 + _source_stream_conv2d_4_source_33_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_buf_3;
  wire _set_flag_489;
  assign _set_flag_489 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_490;
  assign read_rtl_bank_490 = _stream_conv2d_4_source_34_source_ram_raddr;
  reg [1-1:0] _tmp_491;
  assign ram_w16_l512_id8_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17))? _stream_conv2d_4_source_34_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id8_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17))? 1'd1 : 0;
  localparam _tmp_492 = 1;
  wire [_tmp_492-1:0] _tmp_493;
  assign _tmp_493 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17);
  reg [_tmp_492-1:0] __tmp_493_1;
  assign ram_w16_l512_id8_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17))? _stream_conv2d_4_source_34_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id8_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17))? 1'd1 : 0;
  localparam _tmp_494 = 1;
  wire [_tmp_494-1:0] _tmp_495;
  assign _tmp_495 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17);
  reg [_tmp_494-1:0] __tmp_495_1;
  wire signed [16-1:0] read_rtl_rdata_496;
  wire read_rtl_rvalid_497;
  assign read_rtl_rdata_496 = (_tmp_491 == 0)? ram_w16_l512_id8_0_0_rdata : 
                              (_tmp_491 == 1)? ram_w16_l512_id8_1_0_rdata : 0;
  assign read_rtl_rvalid_497 = __tmp_493_1;
  assign _stream_conv2d_4_source_34_source_ram_rdata = (_stream_conv2d_4_source_34_source_sel == 17)? read_rtl_rdata_496 : 'hx;
  reg [16-1:0] __variable_wdata_632;
  assign stream_conv2d_4_source_34_data = __variable_wdata_632;
  reg [32-1:0] _stream_conv2d_4_source_34_source_pat_fsm_16;
  localparam _stream_conv2d_4_source_34_source_pat_fsm_16_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_34_source_pat_all_offset;
  assign _stream_conv2d_4_source_34_source_pat_all_offset = _stream_conv2d_4_source_34_source_offset_buf + _source_stream_conv2d_4_source_34_pat_cur_offset_0 + _source_stream_conv2d_4_source_34_pat_cur_offset_1 + _source_stream_conv2d_4_source_34_pat_cur_offset_2 + _source_stream_conv2d_4_source_34_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_buf_3;
  wire _set_flag_498;
  assign _set_flag_498 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_499;
  assign read_rtl_bank_499 = _stream_conv2d_4_source_35_source_ram_raddr;
  reg [1-1:0] _tmp_500;
  assign ram_w16_l512_id9_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18))? _stream_conv2d_4_source_35_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id9_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18))? 1'd1 : 0;
  localparam _tmp_501 = 1;
  wire [_tmp_501-1:0] _tmp_502;
  assign _tmp_502 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18);
  reg [_tmp_501-1:0] __tmp_502_1;
  assign ram_w16_l512_id9_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18))? _stream_conv2d_4_source_35_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id9_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18))? 1'd1 : 0;
  localparam _tmp_503 = 1;
  wire [_tmp_503-1:0] _tmp_504;
  assign _tmp_504 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18);
  reg [_tmp_503-1:0] __tmp_504_1;
  wire signed [16-1:0] read_rtl_rdata_505;
  wire read_rtl_rvalid_506;
  assign read_rtl_rdata_505 = (_tmp_500 == 0)? ram_w16_l512_id9_0_0_rdata : 
                              (_tmp_500 == 1)? ram_w16_l512_id9_1_0_rdata : 0;
  assign read_rtl_rvalid_506 = __tmp_502_1;
  assign _stream_conv2d_4_source_35_source_ram_rdata = (_stream_conv2d_4_source_35_source_sel == 18)? read_rtl_rdata_505 : 'hx;
  reg [16-1:0] __variable_wdata_633;
  assign stream_conv2d_4_source_35_data = __variable_wdata_633;
  reg [32-1:0] _stream_conv2d_4_source_35_source_pat_fsm_17;
  localparam _stream_conv2d_4_source_35_source_pat_fsm_17_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_35_source_pat_all_offset;
  assign _stream_conv2d_4_source_35_source_pat_all_offset = _stream_conv2d_4_source_35_source_offset_buf + _source_stream_conv2d_4_source_35_pat_cur_offset_0 + _source_stream_conv2d_4_source_35_pat_cur_offset_1 + _source_stream_conv2d_4_source_35_pat_cur_offset_2 + _source_stream_conv2d_4_source_35_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_buf_3;
  wire _set_flag_507;
  assign _set_flag_507 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_508;
  assign read_rtl_bank_508 = _stream_conv2d_4_source_36_source_ram_raddr;
  reg [1-1:0] _tmp_509;
  assign ram_w16_l512_id10_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19))? _stream_conv2d_4_source_36_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id10_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19))? 1'd1 : 0;
  localparam _tmp_510 = 1;
  wire [_tmp_510-1:0] _tmp_511;
  assign _tmp_511 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19);
  reg [_tmp_510-1:0] __tmp_511_1;
  assign ram_w16_l512_id10_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19))? _stream_conv2d_4_source_36_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id10_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19))? 1'd1 : 0;
  localparam _tmp_512 = 1;
  wire [_tmp_512-1:0] _tmp_513;
  assign _tmp_513 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19);
  reg [_tmp_512-1:0] __tmp_513_1;
  wire signed [16-1:0] read_rtl_rdata_514;
  wire read_rtl_rvalid_515;
  assign read_rtl_rdata_514 = (_tmp_509 == 0)? ram_w16_l512_id10_0_0_rdata : 
                              (_tmp_509 == 1)? ram_w16_l512_id10_1_0_rdata : 0;
  assign read_rtl_rvalid_515 = __tmp_511_1;
  assign _stream_conv2d_4_source_36_source_ram_rdata = (_stream_conv2d_4_source_36_source_sel == 19)? read_rtl_rdata_514 : 'hx;
  reg [16-1:0] __variable_wdata_634;
  assign stream_conv2d_4_source_36_data = __variable_wdata_634;
  reg [32-1:0] _stream_conv2d_4_source_36_source_pat_fsm_18;
  localparam _stream_conv2d_4_source_36_source_pat_fsm_18_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_36_source_pat_all_offset;
  assign _stream_conv2d_4_source_36_source_pat_all_offset = _stream_conv2d_4_source_36_source_offset_buf + _source_stream_conv2d_4_source_36_pat_cur_offset_0 + _source_stream_conv2d_4_source_36_pat_cur_offset_1 + _source_stream_conv2d_4_source_36_pat_cur_offset_2 + _source_stream_conv2d_4_source_36_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_buf_3;
  wire _set_flag_516;
  assign _set_flag_516 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_517;
  assign read_rtl_bank_517 = _stream_conv2d_4_source_37_source_ram_raddr;
  reg [1-1:0] _tmp_518;
  assign ram_w16_l512_id11_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20))? _stream_conv2d_4_source_37_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id11_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20))? 1'd1 : 0;
  localparam _tmp_519 = 1;
  wire [_tmp_519-1:0] _tmp_520;
  assign _tmp_520 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20);
  reg [_tmp_519-1:0] __tmp_520_1;
  assign ram_w16_l512_id11_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20))? _stream_conv2d_4_source_37_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id11_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20))? 1'd1 : 0;
  localparam _tmp_521 = 1;
  wire [_tmp_521-1:0] _tmp_522;
  assign _tmp_522 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20);
  reg [_tmp_521-1:0] __tmp_522_1;
  wire signed [16-1:0] read_rtl_rdata_523;
  wire read_rtl_rvalid_524;
  assign read_rtl_rdata_523 = (_tmp_518 == 0)? ram_w16_l512_id11_0_0_rdata : 
                              (_tmp_518 == 1)? ram_w16_l512_id11_1_0_rdata : 0;
  assign read_rtl_rvalid_524 = __tmp_520_1;
  assign _stream_conv2d_4_source_37_source_ram_rdata = (_stream_conv2d_4_source_37_source_sel == 20)? read_rtl_rdata_523 : 'hx;
  reg [16-1:0] __variable_wdata_635;
  assign stream_conv2d_4_source_37_data = __variable_wdata_635;
  reg [32-1:0] _stream_conv2d_4_source_37_source_pat_fsm_19;
  localparam _stream_conv2d_4_source_37_source_pat_fsm_19_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_37_source_pat_all_offset;
  assign _stream_conv2d_4_source_37_source_pat_all_offset = _stream_conv2d_4_source_37_source_offset_buf + _source_stream_conv2d_4_source_37_pat_cur_offset_0 + _source_stream_conv2d_4_source_37_pat_cur_offset_1 + _source_stream_conv2d_4_source_37_pat_cur_offset_2 + _source_stream_conv2d_4_source_37_pat_cur_offset_3;
  wire _set_flag_525;
  assign _set_flag_525 = conv2d_4_comp_fsm == 3;
  reg _tmp_526;
  reg _tmp_527;
  reg _tmp_528;
  reg _tmp_529;
  reg _tmp_530;
  reg _tmp_531;
  reg _tmp_532;
  reg _tmp_533;
  reg _tmp_534;
  reg _tmp_535;
  reg _tmp_536;
  reg _tmp_537;
  reg _tmp_538;
  reg _tmp_539;
  reg _tmp_540;
  reg _tmp_541;
  reg _tmp_542;
  reg _tmp_543;
  reg _tmp_544;
  reg _tmp_545;
  reg _tmp_546;
  reg _tmp_547;
  reg _tmp_548;
  reg _tmp_549;
  reg _tmp_550;
  reg _tmp_551;
  reg _tmp_552;
  reg _tmp_553;
  reg _tmp_554;
  reg _tmp_555;
  reg _tmp_556;
  reg _tmp_557;
  reg _tmp_558;
  localparam _tmp_559 = 33;
  wire [_tmp_559-1:0] _tmp_560;
  assign _tmp_560 = conv2d_4_stream_out_local + conv2d_4_out_page_comp_offset_buf;
  reg [_tmp_559-1:0] _tmp_561;
  reg [_tmp_559-1:0] _tmp_562;
  reg [_tmp_559-1:0] _tmp_563;
  reg [_tmp_559-1:0] _tmp_564;
  reg [_tmp_559-1:0] _tmp_565;
  reg [_tmp_559-1:0] _tmp_566;
  reg [_tmp_559-1:0] _tmp_567;
  reg [_tmp_559-1:0] _tmp_568;
  reg [_tmp_559-1:0] _tmp_569;
  reg [_tmp_559-1:0] _tmp_570;
  reg [_tmp_559-1:0] _tmp_571;
  reg [_tmp_559-1:0] _tmp_572;
  reg [_tmp_559-1:0] _tmp_573;
  reg [_tmp_559-1:0] _tmp_574;
  reg [_tmp_559-1:0] _tmp_575;
  reg [_tmp_559-1:0] _tmp_576;
  reg [_tmp_559-1:0] _tmp_577;
  reg [_tmp_559-1:0] _tmp_578;
  reg [_tmp_559-1:0] _tmp_579;
  reg [_tmp_559-1:0] _tmp_580;
  reg [_tmp_559-1:0] _tmp_581;
  reg [_tmp_559-1:0] _tmp_582;
  reg [_tmp_559-1:0] _tmp_583;
  reg [_tmp_559-1:0] _tmp_584;
  reg [_tmp_559-1:0] _tmp_585;
  reg [_tmp_559-1:0] _tmp_586;
  reg [_tmp_559-1:0] _tmp_587;
  reg [_tmp_559-1:0] _tmp_588;
  reg [_tmp_559-1:0] _tmp_589;
  reg [_tmp_559-1:0] _tmp_590;
  reg [_tmp_559-1:0] _tmp_591;
  reg [_tmp_559-1:0] _tmp_592;
  reg [_tmp_559-1:0] _tmp_593;
  reg [32-1:0] _tmp_594;
  reg [32-1:0] _tmp_595;
  reg [32-1:0] _tmp_596;
  reg [32-1:0] _tmp_597;
  reg [32-1:0] _tmp_598;
  reg [32-1:0] _tmp_599;
  reg [32-1:0] _tmp_600;
  reg [32-1:0] _tmp_601;
  reg [32-1:0] _tmp_602;
  reg [32-1:0] _tmp_603;
  reg [32-1:0] _tmp_604;
  reg [32-1:0] _tmp_605;
  reg [32-1:0] _tmp_606;
  reg [32-1:0] _tmp_607;
  reg [32-1:0] _tmp_608;
  reg [32-1:0] _tmp_609;
  reg [32-1:0] _tmp_610;
  reg [32-1:0] _tmp_611;
  reg [32-1:0] _tmp_612;
  reg [32-1:0] _tmp_613;
  reg [32-1:0] _tmp_614;
  reg [32-1:0] _tmp_615;
  reg [32-1:0] _tmp_616;
  reg [32-1:0] _tmp_617;
  reg [32-1:0] _tmp_618;
  reg [32-1:0] _tmp_619;
  reg [32-1:0] _tmp_620;
  reg [32-1:0] _tmp_621;
  reg [32-1:0] _tmp_622;
  reg [32-1:0] _tmp_623;
  reg [32-1:0] _tmp_624;
  reg [32-1:0] _tmp_625;
  reg [32-1:0] _tmp_626;
  wire [1-1:0] write_rtl_bank_627;
  assign write_rtl_bank_627 = _stream_conv2d_4_sink_50_sink_waddr;
  reg [32-1:0] _stream_conv2d_4_sink_50_sink_fsm_20;
  localparam _stream_conv2d_4_sink_50_sink_fsm_20_init = 0;
  wire _set_flag_628;
  assign _set_flag_628 = conv2d_4_comp_fsm == 4;
  assign _stream_conv2d_4_run_flag = (_set_flag_628)? 1 : 0;
  reg _tmp_629;
  reg _tmp_630;
  reg _tmp_631;
  assign _mul_8_source_stop = _mul_8_stream_oready && 1'd0;
  reg _tmp_632;
  reg _tmp_633;
  reg _tmp_634;
  reg _tmp_635;
  reg _tmp_636;
  reg _tmp_637;
  reg _tmp_638;
  reg _tmp_639;
  reg _tmp_640;
  reg _tmp_641;
  assign _mul_8_sink_start = _tmp_641;
  reg _tmp_642;
  reg _tmp_643;
  reg _tmp_644;
  reg _tmp_645;
  reg _tmp_646;
  reg _tmp_647;
  reg _tmp_648;
  reg _tmp_649;
  reg _tmp_650;
  reg _tmp_651;
  assign _mul_8_sink_stop = _tmp_651;
  reg _tmp_652;
  reg _tmp_653;
  reg _tmp_654;
  reg _tmp_655;
  reg _tmp_656;
  reg _tmp_657;
  reg _tmp_658;
  reg _tmp_659;
  reg _tmp_660;
  reg _tmp_661;
  assign _mul_8_sink_busy = _tmp_661;
  reg _tmp_662;
  assign _mul_8_busy = _mul_8_source_busy || _mul_8_sink_busy || _mul_8_busy_reg;
  reg _tmp_663;
  reg _tmp_664;
  reg _tmp_665;
  assign _mul_9_source_stop = _mul_9_stream_oready && 1'd0;
  reg _tmp_666;
  reg _tmp_667;
  reg _tmp_668;
  reg _tmp_669;
  reg _tmp_670;
  reg _tmp_671;
  reg _tmp_672;
  reg _tmp_673;
  reg _tmp_674;
  reg _tmp_675;
  assign _mul_9_sink_start = _tmp_675;
  reg _tmp_676;
  reg _tmp_677;
  reg _tmp_678;
  reg _tmp_679;
  reg _tmp_680;
  reg _tmp_681;
  reg _tmp_682;
  reg _tmp_683;
  reg _tmp_684;
  reg _tmp_685;
  assign _mul_9_sink_stop = _tmp_685;
  reg _tmp_686;
  reg _tmp_687;
  reg _tmp_688;
  reg _tmp_689;
  reg _tmp_690;
  reg _tmp_691;
  reg _tmp_692;
  reg _tmp_693;
  reg _tmp_694;
  reg _tmp_695;
  assign _mul_9_sink_busy = _tmp_695;
  reg _tmp_696;
  assign _mul_9_busy = _mul_9_source_busy || _mul_9_sink_busy || _mul_9_busy_reg;
  reg _tmp_697;
  reg _tmp_698;
  reg _tmp_699;
  assign _mul_10_source_stop = _mul_10_stream_oready && 1'd0;
  reg _tmp_700;
  reg _tmp_701;
  reg _tmp_702;
  reg _tmp_703;
  reg _tmp_704;
  reg _tmp_705;
  reg _tmp_706;
  reg _tmp_707;
  reg _tmp_708;
  reg _tmp_709;
  assign _mul_10_sink_start = _tmp_709;
  reg _tmp_710;
  reg _tmp_711;
  reg _tmp_712;
  reg _tmp_713;
  reg _tmp_714;
  reg _tmp_715;
  reg _tmp_716;
  reg _tmp_717;
  reg _tmp_718;
  reg _tmp_719;
  assign _mul_10_sink_stop = _tmp_719;
  reg _tmp_720;
  reg _tmp_721;
  reg _tmp_722;
  reg _tmp_723;
  reg _tmp_724;
  reg _tmp_725;
  reg _tmp_726;
  reg _tmp_727;
  reg _tmp_728;
  reg _tmp_729;
  assign _mul_10_sink_busy = _tmp_729;
  reg _tmp_730;
  assign _mul_10_busy = _mul_10_source_busy || _mul_10_sink_busy || _mul_10_busy_reg;
  reg _tmp_731;
  reg _tmp_732;
  reg _tmp_733;
  assign _mul_11_source_stop = _mul_11_stream_oready && 1'd0;
  reg _tmp_734;
  reg _tmp_735;
  reg _tmp_736;
  reg _tmp_737;
  reg _tmp_738;
  reg _tmp_739;
  reg _tmp_740;
  reg _tmp_741;
  reg _tmp_742;
  reg _tmp_743;
  assign _mul_11_sink_start = _tmp_743;
  reg _tmp_744;
  reg _tmp_745;
  reg _tmp_746;
  reg _tmp_747;
  reg _tmp_748;
  reg _tmp_749;
  reg _tmp_750;
  reg _tmp_751;
  reg _tmp_752;
  reg _tmp_753;
  assign _mul_11_sink_stop = _tmp_753;
  reg _tmp_754;
  reg _tmp_755;
  reg _tmp_756;
  reg _tmp_757;
  reg _tmp_758;
  reg _tmp_759;
  reg _tmp_760;
  reg _tmp_761;
  reg _tmp_762;
  reg _tmp_763;
  assign _mul_11_sink_busy = _tmp_763;
  reg _tmp_764;
  assign _mul_11_busy = _mul_11_source_busy || _mul_11_sink_busy || _mul_11_busy_reg;
  reg _tmp_765;
  reg _tmp_766;
  reg _tmp_767;
  assign _mul_12_source_stop = _mul_12_stream_oready && 1'd0;
  reg _tmp_768;
  reg _tmp_769;
  reg _tmp_770;
  reg _tmp_771;
  reg _tmp_772;
  reg _tmp_773;
  reg _tmp_774;
  reg _tmp_775;
  reg _tmp_776;
  reg _tmp_777;
  assign _mul_12_sink_start = _tmp_777;
  reg _tmp_778;
  reg _tmp_779;
  reg _tmp_780;
  reg _tmp_781;
  reg _tmp_782;
  reg _tmp_783;
  reg _tmp_784;
  reg _tmp_785;
  reg _tmp_786;
  reg _tmp_787;
  assign _mul_12_sink_stop = _tmp_787;
  reg _tmp_788;
  reg _tmp_789;
  reg _tmp_790;
  reg _tmp_791;
  reg _tmp_792;
  reg _tmp_793;
  reg _tmp_794;
  reg _tmp_795;
  reg _tmp_796;
  reg _tmp_797;
  assign _mul_12_sink_busy = _tmp_797;
  reg _tmp_798;
  assign _mul_12_busy = _mul_12_source_busy || _mul_12_sink_busy || _mul_12_busy_reg;
  reg _tmp_799;
  reg _tmp_800;
  reg _tmp_801;
  assign _mul_13_source_stop = _mul_13_stream_oready && 1'd0;
  reg _tmp_802;
  reg _tmp_803;
  reg _tmp_804;
  reg _tmp_805;
  reg _tmp_806;
  reg _tmp_807;
  reg _tmp_808;
  reg _tmp_809;
  reg _tmp_810;
  reg _tmp_811;
  assign _mul_13_sink_start = _tmp_811;
  reg _tmp_812;
  reg _tmp_813;
  reg _tmp_814;
  reg _tmp_815;
  reg _tmp_816;
  reg _tmp_817;
  reg _tmp_818;
  reg _tmp_819;
  reg _tmp_820;
  reg _tmp_821;
  assign _mul_13_sink_stop = _tmp_821;
  reg _tmp_822;
  reg _tmp_823;
  reg _tmp_824;
  reg _tmp_825;
  reg _tmp_826;
  reg _tmp_827;
  reg _tmp_828;
  reg _tmp_829;
  reg _tmp_830;
  reg _tmp_831;
  assign _mul_13_sink_busy = _tmp_831;
  reg _tmp_832;
  assign _mul_13_busy = _mul_13_source_busy || _mul_13_sink_busy || _mul_13_busy_reg;
  reg _tmp_833;
  reg _tmp_834;
  reg _tmp_835;
  assign _mul_14_source_stop = _mul_14_stream_oready && 1'd0;
  reg _tmp_836;
  reg _tmp_837;
  reg _tmp_838;
  reg _tmp_839;
  reg _tmp_840;
  reg _tmp_841;
  reg _tmp_842;
  reg _tmp_843;
  reg _tmp_844;
  reg _tmp_845;
  assign _mul_14_sink_start = _tmp_845;
  reg _tmp_846;
  reg _tmp_847;
  reg _tmp_848;
  reg _tmp_849;
  reg _tmp_850;
  reg _tmp_851;
  reg _tmp_852;
  reg _tmp_853;
  reg _tmp_854;
  reg _tmp_855;
  assign _mul_14_sink_stop = _tmp_855;
  reg _tmp_856;
  reg _tmp_857;
  reg _tmp_858;
  reg _tmp_859;
  reg _tmp_860;
  reg _tmp_861;
  reg _tmp_862;
  reg _tmp_863;
  reg _tmp_864;
  reg _tmp_865;
  assign _mul_14_sink_busy = _tmp_865;
  reg _tmp_866;
  assign _mul_14_busy = _mul_14_source_busy || _mul_14_sink_busy || _mul_14_busy_reg;
  reg _tmp_867;
  reg _tmp_868;
  reg _tmp_869;
  assign _mul_15_source_stop = _mul_15_stream_oready && 1'd0;
  reg _tmp_870;
  reg _tmp_871;
  reg _tmp_872;
  reg _tmp_873;
  reg _tmp_874;
  reg _tmp_875;
  reg _tmp_876;
  reg _tmp_877;
  reg _tmp_878;
  reg _tmp_879;
  assign _mul_15_sink_start = _tmp_879;
  reg _tmp_880;
  reg _tmp_881;
  reg _tmp_882;
  reg _tmp_883;
  reg _tmp_884;
  reg _tmp_885;
  reg _tmp_886;
  reg _tmp_887;
  reg _tmp_888;
  reg _tmp_889;
  assign _mul_15_sink_stop = _tmp_889;
  reg _tmp_890;
  reg _tmp_891;
  reg _tmp_892;
  reg _tmp_893;
  reg _tmp_894;
  reg _tmp_895;
  reg _tmp_896;
  reg _tmp_897;
  reg _tmp_898;
  reg _tmp_899;
  assign _mul_15_sink_busy = _tmp_899;
  reg _tmp_900;
  assign _mul_15_busy = _mul_15_source_busy || _mul_15_sink_busy || _mul_15_busy_reg;
  reg _tmp_901;
  reg _tmp_902;
  reg _tmp_903;
  assign _mul_16_source_stop = _mul_16_stream_oready && 1'd0;
  reg _tmp_904;
  reg _tmp_905;
  reg _tmp_906;
  reg _tmp_907;
  reg _tmp_908;
  reg _tmp_909;
  reg _tmp_910;
  reg _tmp_911;
  reg _tmp_912;
  reg _tmp_913;
  assign _mul_16_sink_start = _tmp_913;
  reg _tmp_914;
  reg _tmp_915;
  reg _tmp_916;
  reg _tmp_917;
  reg _tmp_918;
  reg _tmp_919;
  reg _tmp_920;
  reg _tmp_921;
  reg _tmp_922;
  reg _tmp_923;
  assign _mul_16_sink_stop = _tmp_923;
  reg _tmp_924;
  reg _tmp_925;
  reg _tmp_926;
  reg _tmp_927;
  reg _tmp_928;
  reg _tmp_929;
  reg _tmp_930;
  reg _tmp_931;
  reg _tmp_932;
  reg _tmp_933;
  assign _mul_16_sink_busy = _tmp_933;
  reg _tmp_934;
  assign _mul_16_busy = _mul_16_source_busy || _mul_16_sink_busy || _mul_16_busy_reg;
  reg _tmp_935;
  reg _tmp_936;
  reg _tmp_937;
  assign _add_tree_5_source_stop = _add_tree_5_stream_oready && 1'd0;
  reg _tmp_938;
  reg _tmp_939;
  reg _tmp_940;
  reg _tmp_941;
  assign _add_tree_5_sink_start = _tmp_941;
  reg _tmp_942;
  reg _tmp_943;
  reg _tmp_944;
  reg _tmp_945;
  assign _add_tree_5_sink_stop = _tmp_945;
  reg _tmp_946;
  reg _tmp_947;
  reg _tmp_948;
  reg _tmp_949;
  assign _add_tree_5_sink_busy = _tmp_949;
  reg _tmp_950;
  assign _add_tree_5_busy = _add_tree_5_source_busy || _add_tree_5_sink_busy || _add_tree_5_busy_reg;
  reg _tmp_951;
  reg _tmp_952;
  reg _tmp_953;
  reg _tmp_954;
  reg _tmp_955;
  reg _tmp_956;
  reg _tmp_957;
  reg _tmp_958;
  reg _tmp_959;
  reg _tmp_960;
  assign _acc_0_source_stop = _acc_0_stream_oready && 1'd0;
  reg _tmp_961;
  reg _tmp_962;
  reg _tmp_963;
  reg _tmp_964;
  reg _tmp_965;
  reg _tmp_966;
  reg _tmp_967;
  assign _acc_0_sink_start = _tmp_967;
  reg _tmp_968;
  reg _tmp_969;
  reg _tmp_970;
  reg _tmp_971;
  reg _tmp_972;
  reg _tmp_973;
  reg _tmp_974;
  assign _acc_0_sink_stop = _tmp_974;
  reg _tmp_975;
  reg _tmp_976;
  reg _tmp_977;
  reg _tmp_978;
  reg _tmp_979;
  reg _tmp_980;
  reg _tmp_981;
  assign _acc_0_sink_busy = _tmp_981;
  reg _tmp_982;
  assign _acc_0_busy = _acc_0_source_busy || _acc_0_sink_busy || _acc_0_busy_reg;
  reg _tmp_983;
  reg _tmp_984;
  reg _tmp_985;
  assign _mul_rshift_round_clip_6_source_stop = _mul_rshift_round_clip_6_stream_oready && 1'd0;
  reg _tmp_986;
  reg _tmp_987;
  reg _tmp_988;
  reg _tmp_989;
  reg _tmp_990;
  reg _tmp_991;
  reg _tmp_992;
  reg _tmp_993;
  reg _tmp_994;
  reg _tmp_995;
  assign _mul_rshift_round_clip_6_sink_start = _tmp_995;
  reg _tmp_996;
  reg _tmp_997;
  reg _tmp_998;
  reg _tmp_999;
  reg _tmp_1000;
  reg _tmp_1001;
  reg _tmp_1002;
  reg _tmp_1003;
  reg _tmp_1004;
  reg _tmp_1005;
  assign _mul_rshift_round_clip_6_sink_stop = _tmp_1005;
  reg _tmp_1006;
  reg _tmp_1007;
  reg _tmp_1008;
  reg _tmp_1009;
  reg _tmp_1010;
  reg _tmp_1011;
  reg _tmp_1012;
  reg _tmp_1013;
  reg _tmp_1014;
  reg _tmp_1015;
  assign _mul_rshift_round_clip_6_sink_busy = _tmp_1015;
  reg _tmp_1016;
  assign _mul_rshift_round_clip_6_busy = _mul_rshift_round_clip_6_source_busy || _mul_rshift_round_clip_6_sink_busy || _mul_rshift_round_clip_6_busy_reg;
  reg _tmp_1017;
  reg _tmp_1018;
  reg _tmp_1019;
  reg _tmp_1020;
  reg _tmp_1021;
  reg _tmp_1022;
  reg [1-1:0] __variable_wdata_344;
  assign stream_conv2d_4__reduce_reset_data = __variable_wdata_344;
  reg _tmp_1023;
  reg _tmp_1024;
  reg _tmp_1025;
  reg _tmp_1026;
  assign _stream_conv2d_4_source_stop = _stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3));
  localparam _tmp_1027 = 1;
  wire [_tmp_1027-1:0] _tmp_1028;
  assign _tmp_1028 = _stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3);
  reg [_tmp_1027-1:0] _tmp_1029;
  localparam _tmp_1030 = 1;
  wire [_tmp_1030-1:0] _tmp_1031;
  assign _tmp_1031 = _stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3);
  reg [_tmp_1030-1:0] _tmp_1032;
  reg _tmp_1033;
  reg _tmp_1034;
  reg _tmp_1035;
  reg _tmp_1036;
  reg _tmp_1037;
  reg _tmp_1038;
  reg _tmp_1039;
  reg _tmp_1040;
  reg _tmp_1041;
  reg _tmp_1042;
  reg _tmp_1043;
  reg _tmp_1044;
  reg _tmp_1045;
  reg _tmp_1046;
  reg _tmp_1047;
  reg _tmp_1048;
  reg _tmp_1049;
  reg _tmp_1050;
  reg _tmp_1051;
  reg _tmp_1052;
  reg _tmp_1053;
  reg _tmp_1054;
  reg _tmp_1055;
  reg _tmp_1056;
  reg _tmp_1057;
  reg _tmp_1058;
  reg _tmp_1059;
  reg _tmp_1060;
  reg _tmp_1061;
  reg _tmp_1062;
  reg _tmp_1063;
  reg _tmp_1064;
  reg _tmp_1065;
  assign _stream_conv2d_4_sink_start = _tmp_1065;
  reg _tmp_1066;
  reg _tmp_1067;
  reg _tmp_1068;
  reg _tmp_1069;
  reg _tmp_1070;
  reg _tmp_1071;
  reg _tmp_1072;
  reg _tmp_1073;
  reg _tmp_1074;
  reg _tmp_1075;
  reg _tmp_1076;
  reg _tmp_1077;
  reg _tmp_1078;
  reg _tmp_1079;
  reg _tmp_1080;
  reg _tmp_1081;
  reg _tmp_1082;
  reg _tmp_1083;
  reg _tmp_1084;
  reg _tmp_1085;
  reg _tmp_1086;
  reg _tmp_1087;
  reg _tmp_1088;
  reg _tmp_1089;
  reg _tmp_1090;
  reg _tmp_1091;
  reg _tmp_1092;
  reg _tmp_1093;
  reg _tmp_1094;
  reg _tmp_1095;
  reg _tmp_1096;
  reg _tmp_1097;
  reg _tmp_1098;
  assign _stream_conv2d_4_sink_stop = _tmp_1098;
  reg _tmp_1099;
  reg _tmp_1100;
  reg _tmp_1101;
  reg _tmp_1102;
  reg _tmp_1103;
  reg _tmp_1104;
  reg _tmp_1105;
  reg _tmp_1106;
  reg _tmp_1107;
  reg _tmp_1108;
  reg _tmp_1109;
  reg _tmp_1110;
  reg _tmp_1111;
  reg _tmp_1112;
  reg _tmp_1113;
  reg _tmp_1114;
  reg _tmp_1115;
  reg _tmp_1116;
  reg _tmp_1117;
  reg _tmp_1118;
  reg _tmp_1119;
  reg _tmp_1120;
  reg _tmp_1121;
  reg _tmp_1122;
  reg _tmp_1123;
  reg _tmp_1124;
  reg _tmp_1125;
  reg _tmp_1126;
  reg _tmp_1127;
  reg _tmp_1128;
  reg _tmp_1129;
  reg _tmp_1130;
  reg _tmp_1131;
  assign _stream_conv2d_4_sink_busy = _tmp_1131;
  reg _tmp_1132;
  assign _stream_conv2d_4_busy = _stream_conv2d_4_source_busy || _stream_conv2d_4_sink_busy || _stream_conv2d_4_busy_reg;
  wire conv2d_4_dma_out_mask_0;
  assign conv2d_4_dma_out_mask_0 = conv2d_4_out_row_count + 0 >= cparam_conv2d_4_out_num_row;
  wire [32-1:0] _dma_write_packed_high_local_size_1133;
  assign _dma_write_packed_high_local_size_1133 = conv2d_4_next_out_write_size >> 1;
  wire [1-1:0] _dma_write_packed_low_local_size_1134;
  assign _dma_write_packed_low_local_size_1134 = conv2d_4_next_out_write_size & { 1{ 1'd1 } };
  wire [32-1:0] _dma_write_packed_local_packed_size_1135;
  assign _dma_write_packed_local_packed_size_1135 = (_dma_write_packed_low_local_size_1134 > 0)? _dma_write_packed_high_local_size_1133 + 1 : _dma_write_packed_high_local_size_1133;
  wire [32-1:0] mask_addr_shifted_1136;
  assign mask_addr_shifted_1136 = conv2d_4_objaddr + (conv2d_4_out_base_offset + cparam_conv2d_4_out_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1137;
  assign mask_addr_masked_1137 = mask_addr_shifted_1136 << 2;
  reg [32-1:0] _maxi_write_req_fsm;
  localparam _maxi_write_req_fsm_init = 0;
  reg [33-1:0] _maxi_write_cur_global_size;
  reg _maxi_write_cont;
  wire [8-1:0] pack_write_req_op_sel_1138;
  wire [32-1:0] pack_write_req_local_addr_1139;
  wire [32-1:0] pack_write_req_local_stride_1140;
  wire [33-1:0] pack_write_req_size_1141;
  wire [32-1:0] pack_write_req_local_blocksize_1142;
  assign pack_write_req_op_sel_1138 = _maxi_write_op_sel;
  assign pack_write_req_local_addr_1139 = _maxi_write_local_addr;
  assign pack_write_req_local_stride_1140 = _maxi_write_local_stride;
  assign pack_write_req_size_1141 = _maxi_write_local_size;
  assign pack_write_req_local_blocksize_1142 = _maxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_1143;
  assign pack_write_req_packed_1143 = { pack_write_req_op_sel_1138, pack_write_req_local_addr_1139, pack_write_req_local_stride_1140, pack_write_req_size_1141, pack_write_req_local_blocksize_1142 };
  localparam _tmp_1144 = 1;
  wire [_tmp_1144-1:0] _tmp_1145;
  assign _tmp_1145 = !_maxi_write_req_fifo_almost_full;
  reg [_tmp_1144-1:0] __tmp_1145_1;
  wire [32-1:0] mask_addr_shifted_1146;
  assign mask_addr_shifted_1146 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1147;
  assign mask_addr_masked_1147 = mask_addr_shifted_1146 << 2;
  wire [32-1:0] mask_addr_shifted_1148;
  assign mask_addr_shifted_1148 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1149;
  assign mask_addr_masked_1149 = mask_addr_shifted_1148 << 2;
  wire [32-1:0] mask_addr_shifted_1150;
  assign mask_addr_shifted_1150 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1151;
  assign mask_addr_masked_1151 = mask_addr_shifted_1150 << 2;
  wire [32-1:0] mask_addr_shifted_1152;
  assign mask_addr_shifted_1152 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1153;
  assign mask_addr_masked_1153 = mask_addr_shifted_1152 << 2;
  wire [32-1:0] mask_addr_shifted_1154;
  assign mask_addr_shifted_1154 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1155;
  assign mask_addr_masked_1155 = mask_addr_shifted_1154 << 2;
  wire [32-1:0] mask_addr_shifted_1156;
  assign mask_addr_shifted_1156 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1157;
  assign mask_addr_masked_1157 = mask_addr_shifted_1156 << 2;
  wire [8-1:0] pack_write_req_op_sel_1158;
  wire [32-1:0] pack_write_req_local_addr_1159;
  wire [32-1:0] pack_write_req_local_stride_1160;
  wire [33-1:0] pack_write_req_size_1161;
  wire [32-1:0] pack_write_req_local_blocksize_1162;
  assign pack_write_req_op_sel_1158 = _maxi_write_op_sel;
  assign pack_write_req_local_addr_1159 = _maxi_write_local_addr;
  assign pack_write_req_local_stride_1160 = _maxi_write_local_stride;
  assign pack_write_req_size_1161 = _maxi_write_cur_global_size;
  assign pack_write_req_local_blocksize_1162 = _maxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_1163;
  assign pack_write_req_packed_1163 = { pack_write_req_op_sel_1158, pack_write_req_local_addr_1159, pack_write_req_local_stride_1160, pack_write_req_size_1161, pack_write_req_local_blocksize_1162 };
  assign _maxi_write_req_fifo_wdata = ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))? pack_write_req_packed_1163 : 
                                      ((_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full)? pack_write_req_packed_1143 : 'hx;
  assign _maxi_write_req_fifo_enq = ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))? (_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6) && !_maxi_write_req_fifo_almost_full : 
                                    ((_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full)? (_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full && !_maxi_write_req_fifo_almost_full : 0;
  localparam _tmp_1164 = 1;
  wire [_tmp_1164-1:0] _tmp_1165;
  assign _tmp_1165 = !_maxi_write_req_fifo_almost_full;
  reg [_tmp_1164-1:0] __tmp_1165_1;
  reg _maxi_waddr_cond_0_1;
  reg [32-1:0] _maxi_write_data_fsm;
  localparam _maxi_write_data_fsm_init = 0;
  reg [32-1:0] read_burst_packed_fsm_24;
  localparam read_burst_packed_fsm_24_init = 0;
  reg [9-1:0] read_burst_packed_addr_1166;
  reg [9-1:0] read_burst_packed_stride_1167;
  reg [33-1:0] read_burst_packed_length_1168;
  reg read_burst_packed_rvalid_1169;
  reg read_burst_packed_rlast_1170;
  wire [8-1:0] read_burst_packed_ram_addr_1171;
  assign read_burst_packed_ram_addr_1171 = read_burst_packed_addr_1166 >> 1;
  assign ram_w16_l512_id0_0_1_addr = ((read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1169 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1171 : 'hx;
  assign ram_w16_l512_id0_0_1_enable = ((read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1169 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  localparam _tmp_1172 = 1;
  wire [_tmp_1172-1:0] _tmp_1173;
  assign _tmp_1173 = (read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1169 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1172-1:0] __tmp_1173_1;
  wire [16-1:0] read_burst_packed_ram_rdata_1174;
  assign read_burst_packed_ram_rdata_1174 = ram_w16_l512_id0_0_1_rdata;
  wire [8-1:0] read_burst_packed_ram_addr_1175;
  assign read_burst_packed_ram_addr_1175 = read_burst_packed_addr_1166 >> 1;
  assign ram_w16_l512_id0_1_1_addr = ((read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1169 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1175 : 'hx;
  assign ram_w16_l512_id0_1_1_enable = ((read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1169 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  localparam _tmp_1176 = 1;
  wire [_tmp_1176-1:0] _tmp_1177;
  assign _tmp_1177 = (read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1169 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1176-1:0] __tmp_1177_1;
  wire [16-1:0] read_burst_packed_ram_rdata_1178;
  assign read_burst_packed_ram_rdata_1178 = ram_w16_l512_id0_1_1_rdata;
  wire [32-1:0] read_burst_packed_rdata_1179;
  assign read_burst_packed_rdata_1179 = { read_burst_packed_ram_rdata_1178, read_burst_packed_ram_rdata_1174 };
  reg _maxi_wdata_cond_0_1;
  wire conv2d_4_update_filter;
  assign conv2d_4_update_filter = (cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) || (cparam_conv2d_4_data_stationary == 1) && !cparam_conv2d_4_keep_filter;
  wire conv2d_4_update_act;
  assign conv2d_4_update_act = (cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count) || (cparam_conv2d_4_data_stationary == 0);
  wire conv2d_4_mux_next_dma_flag_0;
  assign conv2d_4_mux_next_dma_flag_0 = (conv2d_4_row_select == 0)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_0 : 
                                        (conv2d_4_row_select == 1)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_2 : 
                                        (conv2d_4_row_select == 2)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_1 : 1'd0;
  wire conv2d_4_mux_next_dma_flag_1;
  assign conv2d_4_mux_next_dma_flag_1 = (conv2d_4_row_select == 0)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_1 : 
                                        (conv2d_4_row_select == 1)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_0 : 
                                        (conv2d_4_row_select == 2)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_2 : 1'd0;
  wire conv2d_4_mux_next_dma_flag_2;
  assign conv2d_4_mux_next_dma_flag_2 = (conv2d_4_row_select == 0)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_2 : 
                                        (conv2d_4_row_select == 1)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_1 : 
                                        (conv2d_4_row_select == 2)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_0 : 1'd0;
  reg [32-1:0] max_pool_serial_6_objaddr;
  reg [32-1:0] max_pool_serial_6_arg_objaddr_0;
  reg [32-1:0] control_max_pool_serial_6;
  localparam control_max_pool_serial_6_init = 0;
  reg _control_max_pool_serial_6_called;
  wire signed [32-1:0] max_pool_serial_6_act_base_offset;
  reg signed [32-1:0] max_pool_serial_6_act_base_offset_row;
  reg signed [32-1:0] max_pool_serial_6_act_base_offset_bat;
  assign max_pool_serial_6_act_base_offset = max_pool_serial_6_act_base_offset_row + max_pool_serial_6_act_base_offset_bat;
  wire signed [32-1:0] max_pool_serial_6_out_base_offset;
  reg signed [32-1:0] max_pool_serial_6_out_base_offset_row;
  reg signed [32-1:0] max_pool_serial_6_out_base_offset_bat;
  assign max_pool_serial_6_out_base_offset = max_pool_serial_6_out_base_offset_row + max_pool_serial_6_out_base_offset_bat;
  reg [32-1:0] max_pool_serial_6_col_count;
  reg [32-1:0] max_pool_serial_6_row_count;
  reg [32-1:0] max_pool_serial_6_bat_count;
  reg [32-1:0] max_pool_serial_6_prev_row_count;
  reg [32-1:0] max_pool_serial_6_prev_bat_count;
  reg [32-1:0] max_pool_serial_6_stream_act_local;
  reg [32-1:0] max_pool_serial_6_stream_out_local;
  reg max_pool_serial_6_act_page;
  reg [32-1:0] max_pool_serial_6_act_page_comp_offset;
  reg [32-1:0] max_pool_serial_6_act_page_dma_offset;
  reg max_pool_serial_6_out_page;
  reg [32-1:0] max_pool_serial_6_out_page_comp_offset;
  reg [32-1:0] max_pool_serial_6_out_page_dma_offset;
  reg max_pool_serial_6_skip_read_act;
  reg max_pool_serial_6_skip_comp;
  reg max_pool_serial_6_skip_write_out;
  reg [32-1:0] max_pool_serial_6_comp_count;
  reg [32-1:0] max_pool_serial_6_out_count;
  wire max_pool_serial_6_dma_pad_mask_0;
  assign max_pool_serial_6_dma_pad_mask_0 = (max_pool_serial_6_row_count + 0 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count + 0 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire max_pool_serial_6_dma_pad_mask_1;
  assign max_pool_serial_6_dma_pad_mask_1 = (max_pool_serial_6_row_count + 1 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count + 1 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire [32-1:0] mask_addr_shifted_1180;
  assign mask_addr_shifted_1180 = max_pool_serial_6_arg_objaddr_0 + (max_pool_serial_6_act_base_offset + cparam_max_pool_serial_6_act_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1181;
  assign mask_addr_masked_1181 = mask_addr_shifted_1180 << 2;
  reg [32-1:0] write_burst_fsm_25;
  localparam write_burst_fsm_25_init = 0;
  reg [12-1:0] write_burst_addr_1182;
  reg [12-1:0] write_burst_stride_1183;
  reg [33-1:0] write_burst_length_1184;
  reg write_burst_done_1185;
  assign ram_w32_l4096_id0_1_addr = ((write_burst_fsm_25 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_1182 : 'hx;
  assign ram_w32_l4096_id0_1_wdata = ((write_burst_fsm_25 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l4096_id0_1_wenable = ((write_burst_fsm_25 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l4096_id0_1_enable = ((write_burst_fsm_25 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [32-1:0] mask_addr_shifted_1186;
  assign mask_addr_shifted_1186 = max_pool_serial_6_arg_objaddr_0 + (max_pool_serial_6_act_base_offset + cparam_max_pool_serial_6_act_offset_values_1) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1187;
  assign mask_addr_masked_1187 = mask_addr_shifted_1186 << 2;
  reg [32-1:0] max_pool_serial_6_comp_fsm;
  localparam max_pool_serial_6_comp_fsm_init = 0;
  reg [32-1:0] max_pool_serial_6_act_page_comp_offset_buf;
  reg [32-1:0] max_pool_serial_6_out_page_comp_offset_buf;
  reg [32-1:0] max_pool_serial_6_row_count_buf;
  wire max_pool_serial_6_stream_pad_mask_0_0;
  assign max_pool_serial_6_stream_pad_mask_0_0 = (max_pool_serial_6_col_count + 0 < cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_col_count + 0 >= cparam_max_pool_serial_6_act_num_col + cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_row_count_buf + 0 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count_buf + 0 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire max_pool_serial_6_stream_pad_mask_0_1;
  assign max_pool_serial_6_stream_pad_mask_0_1 = (max_pool_serial_6_col_count + 1 < cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_col_count + 1 >= cparam_max_pool_serial_6_act_num_col + cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_row_count_buf + 0 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count_buf + 0 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire max_pool_serial_6_stream_pad_mask_1_0;
  assign max_pool_serial_6_stream_pad_mask_1_0 = (max_pool_serial_6_col_count + 0 < cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_col_count + 0 >= cparam_max_pool_serial_6_act_num_col + cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_row_count_buf + 1 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count_buf + 1 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire max_pool_serial_6_stream_pad_mask_1_1;
  assign max_pool_serial_6_stream_pad_mask_1_1 = (max_pool_serial_6_col_count + 1 < cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_col_count + 1 >= cparam_max_pool_serial_6_act_num_col + cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_row_count_buf + 1 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count_buf + 1 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  reg [4-1:0] max_pool_serial_6_stream_pad_masks;
  wire [3-1:0] stream_max_pool_serial_6_parameter_0_data;
  wire [32-1:0] stream_max_pool_serial_6_source_1_data;
  wire [4-1:0] stream_max_pool_serial_6_parameter_2_data;
  wire [1-1:0] stream_max_pool_serial_6__reduce_reset_data;
  reg __stream_max_pool_serial_6_stream_ivalid_1;
  reg __stream_max_pool_serial_6_stream_ivalid_2;
  reg __stream_max_pool_serial_6_stream_ivalid_3;
  reg __stream_max_pool_serial_6_stream_ivalid_4;
  reg __stream_max_pool_serial_6_stream_ivalid_5;
  reg [32-1:0] _counter_data_932;
  reg [32-1:0] _counter_count_932;
  wire _counter_reset_cond_932;
  assign _counter_reset_cond_932 = stream_max_pool_serial_6__reduce_reset_data;
  wire [32-1:0] _counter_current_count_932;
  assign _counter_current_count_932 = (_counter_reset_cond_932)? 1'sd0 : _counter_count_932;
  wire [16-1:0] _slice_data_938;
  assign _slice_data_938 = stream_max_pool_serial_6_source_1_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_939;
  assign _reinterpretcast_src_939 = _slice_data_938;
  wire signed [16-1:0] _reinterpretcast_data_939;
  assign _reinterpretcast_data_939 = _reinterpretcast_src_939;
  wire [16-1:0] _slice_data_942;
  assign _slice_data_942 = stream_max_pool_serial_6_source_1_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_943;
  assign _reinterpretcast_src_943 = _slice_data_942;
  wire signed [16-1:0] _reinterpretcast_data_943;
  assign _reinterpretcast_data_943 = _reinterpretcast_src_943;
  reg [4-1:0] __delay_data_1390__variable_930;
  reg signed [16-1:0] __delay_data_1391_reinterpretcast_939;
  reg [1-1:0] __delay_data_1393__variable_931;
  reg [3-1:0] __delay_data_1396__variable_928;
  reg signed [16-1:0] __delay_data_1399_reinterpretcast_943;
  reg [1-1:0] _pointer_data_935;
  reg signed [16-1:0] __delay_data_1392__delay_1391_reinterpretcast_939;
  reg [1-1:0] __delay_data_1394__delay_1393__variable_931;
  reg [3-1:0] __delay_data_1397__delay_1396__variable_928;
  reg signed [16-1:0] __delay_data_1400__delay_1399_reinterpretcast_943;
  reg signed [17-1:0] _cond_data_945;
  reg signed [17-1:0] _cond_data_950;
  reg [1-1:0] __delay_data_1395__delay_1394__delay_1393__variable_931;
  reg [3-1:0] __delay_data_1398__delay_1397__delay_1396__variable_928;
  reg [1-1:0] __variable_wdata_327;
  assign _reduce_max_17__reduce_reset_data = __variable_wdata_327;
  reg signed [16-1:0] __variable_wdata_325;
  assign _reduce_max_17_x_data = __variable_wdata_325;
  reg [32-1:0] __variable_wdata_326;
  assign _reduce_max_17_size_data = __variable_wdata_326;
  assign __reduce_max_17_is_root = ((_stream_max_pool_serial_6_busy)? 0 : 1) && 1;
  assign __reduce_max_17_stream_oready = ((_stream_max_pool_serial_6_busy)? _stream_max_pool_serial_6_stream_oready : 1) && __reduce_max_17_stream_internal_oready;
  reg [1-1:0] __variable_wdata_334;
  assign _reduce_max_18__reduce_reset_data = __variable_wdata_334;
  reg signed [16-1:0] __variable_wdata_332;
  assign _reduce_max_18_x_data = __variable_wdata_332;
  reg [32-1:0] __variable_wdata_333;
  assign _reduce_max_18_size_data = __variable_wdata_333;
  assign __reduce_max_18_is_root = ((_stream_max_pool_serial_6_busy)? 0 : 1) && 1;
  assign __reduce_max_18_stream_oready = ((_stream_max_pool_serial_6_busy)? _stream_max_pool_serial_6_stream_oready : 1) && __reduce_max_18_stream_internal_oready;
  assign _stream_max_pool_serial_6_stream_internal_oready = ((_stream_max_pool_serial_6_busy)? __reduce_max_18_stream_internal_oready : 1) && (((_stream_max_pool_serial_6_busy)? __reduce_max_17_stream_internal_oready : 1) && 1);
  wire signed [16-1:0] __substreamoutput_data_947;
  assign __substreamoutput_data_947 = _reduce_max_17_data_data;
  wire [1-1:0] __substreamoutput_data_948;
  assign __substreamoutput_data_948 = _reduce_max_17_valid_data;
  wire signed [16-1:0] _reinterpretcast_src_949;
  assign _reinterpretcast_src_949 = __substreamoutput_data_947;
  wire signed [16-1:0] _reinterpretcast_data_949;
  assign _reinterpretcast_data_949 = _reinterpretcast_src_949;
  wire signed [16-1:0] __substreamoutput_data_952;
  assign __substreamoutput_data_952 = _reduce_max_18_data_data;
  wire signed [16-1:0] _reinterpretcast_src_954;
  assign _reinterpretcast_src_954 = __substreamoutput_data_952;
  wire signed [16-1:0] _reinterpretcast_data_954;
  assign _reinterpretcast_data_954 = _reinterpretcast_src_954;
  wire [32-1:0] _cat_data_955;
  assign _cat_data_955 = { _reinterpretcast_data_954, _reinterpretcast_data_949 };
  wire [1-1:0] stream_max_pool_serial_6_sink_7_data;
  assign stream_max_pool_serial_6_sink_7_data = __substreamoutput_data_948;
  wire [32-1:0] stream_max_pool_serial_6_sink_6_data;
  assign stream_max_pool_serial_6_sink_6_data = _cat_data_955;
  wire _set_flag_1188;
  assign _set_flag_1188 = max_pool_serial_6_comp_fsm == 4;
  reg [3-1:0] __variable_wdata_928;
  assign stream_max_pool_serial_6_parameter_0_data = __variable_wdata_928;
  wire _set_flag_1189;
  assign _set_flag_1189 = max_pool_serial_6_comp_fsm == 4;
  reg [4-1:0] __variable_wdata_930;
  assign stream_max_pool_serial_6_parameter_2_data = __variable_wdata_930;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_0;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_1;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_2;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_3;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_0;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_1;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_2;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_3;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_count_0;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_count_1;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_count_2;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_count_3;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_buf_0;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_buf_1;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_buf_2;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_buf_3;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_buf_0;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_buf_1;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_buf_2;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_buf_3;
  wire _set_flag_1190;
  assign _set_flag_1190 = max_pool_serial_6_comp_fsm == 4;
  assign ram_w32_l4096_id0_0_addr = (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_1_source_ram_renable && (_stream_max_pool_serial_6_source_1_source_sel == 1))? _stream_max_pool_serial_6_source_1_source_ram_raddr : 'hx;
  assign ram_w32_l4096_id0_0_enable = (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_1_source_ram_renable && (_stream_max_pool_serial_6_source_1_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_1191 = 1;
  wire [_tmp_1191-1:0] _tmp_1192;
  assign _tmp_1192 = _stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_1_source_ram_renable && (_stream_max_pool_serial_6_source_1_source_sel == 1);
  reg [_tmp_1191-1:0] __tmp_1192_1;
  assign _stream_max_pool_serial_6_source_1_source_ram_rdata = (_stream_max_pool_serial_6_source_1_source_sel == 1)? ram_w32_l4096_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_929;
  assign stream_max_pool_serial_6_source_1_data = __variable_wdata_929;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_pat_fsm_0;
  localparam _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_max_pool_serial_6_source_1_source_pat_all_offset;
  assign _stream_max_pool_serial_6_source_1_source_pat_all_offset = _stream_max_pool_serial_6_source_1_source_offset_buf + _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 + _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 + _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 + _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3;
  wire _set_flag_1193;
  assign _set_flag_1193 = max_pool_serial_6_comp_fsm == 4;
  reg _tmp_1194;
  reg _tmp_1195;
  reg _tmp_1196;
  reg _tmp_1197;
  reg _tmp_1198;
  reg _tmp_1199;
  reg _tmp_1200;
  localparam _tmp_1201 = 33;
  wire [_tmp_1201-1:0] _tmp_1202;
  assign _tmp_1202 = max_pool_serial_6_stream_out_local + max_pool_serial_6_out_page_comp_offset_buf;
  reg [_tmp_1201-1:0] _tmp_1203;
  reg [_tmp_1201-1:0] _tmp_1204;
  reg [_tmp_1201-1:0] _tmp_1205;
  reg [_tmp_1201-1:0] _tmp_1206;
  reg [_tmp_1201-1:0] _tmp_1207;
  reg [_tmp_1201-1:0] _tmp_1208;
  reg [_tmp_1201-1:0] _tmp_1209;
  reg [8-1:0] _tmp_1210;
  reg [8-1:0] _tmp_1211;
  reg [8-1:0] _tmp_1212;
  reg [8-1:0] _tmp_1213;
  reg [8-1:0] _tmp_1214;
  reg [8-1:0] _tmp_1215;
  reg [8-1:0] _tmp_1216;
  assign ram_w32_l1024_id0_0_wdata = (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_6_sink_wenable && (_stream_max_pool_serial_6_sink_6_sink_sel == 2))? _stream_max_pool_serial_6_sink_6_sink_wdata : 'hx;
  assign ram_w32_l1024_id0_0_wenable = (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_6_sink_wenable && (_stream_max_pool_serial_6_sink_6_sink_sel == 2))? 1'd1 : 0;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_fsm_1;
  localparam _stream_max_pool_serial_6_sink_6_sink_fsm_1_init = 0;
  wire _set_flag_1217;
  assign _set_flag_1217 = max_pool_serial_6_comp_fsm == 5;
  assign _stream_max_pool_serial_6_run_flag = (_set_flag_1217)? 1 : 0;
  reg _tmp_1218;
  reg _tmp_1219;
  reg _tmp_1220;
  reg _tmp_1221;
  reg _tmp_1222;
  reg _tmp_1223;
  reg _tmp_1224;
  reg _tmp_1225;
  reg _tmp_1226;
  reg _tmp_1227;
  assign __reduce_max_17_source_stop = __reduce_max_17_stream_oready && 1'd0;
  reg _tmp_1228;
  reg _tmp_1229;
  reg _tmp_1230;
  assign __reduce_max_17_sink_start = _tmp_1230;
  reg _tmp_1231;
  reg _tmp_1232;
  reg _tmp_1233;
  assign __reduce_max_17_sink_stop = _tmp_1233;
  reg _tmp_1234;
  reg _tmp_1235;
  reg _tmp_1236;
  assign __reduce_max_17_sink_busy = _tmp_1236;
  reg _tmp_1237;
  assign __reduce_max_17_busy = __reduce_max_17_source_busy || __reduce_max_17_sink_busy || __reduce_max_17_busy_reg;
  reg _tmp_1238;
  reg _tmp_1239;
  reg _tmp_1240;
  reg _tmp_1241;
  reg _tmp_1242;
  reg _tmp_1243;
  reg _tmp_1244;
  reg _tmp_1245;
  reg _tmp_1246;
  reg _tmp_1247;
  assign __reduce_max_18_source_stop = __reduce_max_18_stream_oready && 1'd0;
  reg _tmp_1248;
  reg _tmp_1249;
  reg _tmp_1250;
  assign __reduce_max_18_sink_start = _tmp_1250;
  reg _tmp_1251;
  reg _tmp_1252;
  reg _tmp_1253;
  assign __reduce_max_18_sink_stop = _tmp_1253;
  reg _tmp_1254;
  reg _tmp_1255;
  reg _tmp_1256;
  assign __reduce_max_18_sink_busy = _tmp_1256;
  reg _tmp_1257;
  assign __reduce_max_18_busy = __reduce_max_18_source_busy || __reduce_max_18_sink_busy || __reduce_max_18_busy_reg;
  reg _tmp_1258;
  reg _tmp_1259;
  reg _tmp_1260;
  reg _tmp_1261;
  reg _tmp_1262;
  reg _tmp_1263;
  reg [1-1:0] __variable_wdata_931;
  assign stream_max_pool_serial_6__reduce_reset_data = __variable_wdata_931;
  reg _tmp_1264;
  reg _tmp_1265;
  reg _tmp_1266;
  reg _tmp_1267;
  assign _stream_max_pool_serial_6_source_stop = _stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3));
  localparam _tmp_1268 = 1;
  wire [_tmp_1268-1:0] _tmp_1269;
  assign _tmp_1269 = _stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3);
  reg [_tmp_1268-1:0] _tmp_1270;
  localparam _tmp_1271 = 1;
  wire [_tmp_1271-1:0] _tmp_1272;
  assign _tmp_1272 = _stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3);
  reg [_tmp_1271-1:0] _tmp_1273;
  reg _tmp_1274;
  reg _tmp_1275;
  reg _tmp_1276;
  reg _tmp_1277;
  reg _tmp_1278;
  reg _tmp_1279;
  reg _tmp_1280;
  assign _stream_max_pool_serial_6_sink_start = _tmp_1280;
  reg _tmp_1281;
  reg _tmp_1282;
  reg _tmp_1283;
  reg _tmp_1284;
  reg _tmp_1285;
  reg _tmp_1286;
  reg _tmp_1287;
  assign _stream_max_pool_serial_6_sink_stop = _tmp_1287;
  reg _tmp_1288;
  reg _tmp_1289;
  reg _tmp_1290;
  reg _tmp_1291;
  reg _tmp_1292;
  reg _tmp_1293;
  reg _tmp_1294;
  assign _stream_max_pool_serial_6_sink_busy = _tmp_1294;
  reg _tmp_1295;
  assign _stream_max_pool_serial_6_busy = _stream_max_pool_serial_6_source_busy || _stream_max_pool_serial_6_sink_busy || _stream_max_pool_serial_6_busy_reg;
  wire [32-1:0] mask_addr_shifted_1296;
  assign mask_addr_shifted_1296 = max_pool_serial_6_objaddr + max_pool_serial_6_out_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1297;
  assign mask_addr_masked_1297 = mask_addr_shifted_1296 << 2;
  reg [32-1:0] read_burst_fsm_26;
  localparam read_burst_fsm_26_init = 0;
  reg [10-1:0] read_burst_addr_1298;
  reg [10-1:0] read_burst_stride_1299;
  reg [33-1:0] read_burst_length_1300;
  reg read_burst_rvalid_1301;
  reg read_burst_rlast_1302;
  localparam _tmp_1303 = 1;
  wire [_tmp_1303-1:0] _tmp_1304;
  assign _tmp_1304 = (read_burst_fsm_26 == 1) && (!read_burst_rvalid_1301 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1303-1:0] __tmp_1304_1;
  wire [32-1:0] read_burst_rdata_1305;
  assign read_burst_rdata_1305 = ram_w32_l1024_id0_1_rdata;
  reg _maxi_wdata_cond_1_1;
  reg [32-1:0] matmul_23_objaddr;
  reg [32-1:0] matmul_23_arg_objaddr_0;
  reg [32-1:0] matmul_23_arg_objaddr_1;
  reg [32-1:0] matmul_23_arg_objaddr_2;
  reg [32-1:0] matmul_23_arg_objaddr_3;
  reg [32-1:0] control_matmul_23;
  localparam control_matmul_23_init = 0;
  reg _control_matmul_23_called;
  wire signed [32-1:0] matmul_23_act_base_offset;
  reg signed [32-1:0] matmul_23_act_base_offset_row;
  reg signed [32-1:0] matmul_23_act_base_offset_bat;
  assign matmul_23_act_base_offset = matmul_23_act_base_offset_row + matmul_23_act_base_offset_bat;
  reg signed [32-1:0] matmul_23_filter_base_offset;
  reg [32-1:0] matmul_23_next_stream_num_ops;
  wire signed [32-1:0] matmul_23_out_base_offset;
  reg signed [32-1:0] matmul_23_out_base_offset_val;
  reg signed [32-1:0] matmul_23_out_base_offset_col;
  reg signed [32-1:0] matmul_23_out_base_offset_row;
  reg signed [32-1:0] matmul_23_out_base_offset_bat;
  reg signed [32-1:0] matmul_23_out_base_offset_och;
  assign matmul_23_out_base_offset = matmul_23_out_base_offset_val + matmul_23_out_base_offset_col + matmul_23_out_base_offset_row + matmul_23_out_base_offset_bat + matmul_23_out_base_offset_och;
  reg matmul_23_dma_flag_0;
  reg [32-1:0] matmul_23_sync_comp_count;
  reg [32-1:0] matmul_23_sync_out_count;
  reg [32-1:0] matmul_23_write_count;
  reg [32-1:0] matmul_23_next_out_write_size;
  reg [32-1:0] matmul_23_col_count;
  reg [32-1:0] matmul_23_row_count;
  reg [32-1:0] matmul_23_bat_count;
  reg [32-1:0] matmul_23_och_count;
  reg [1-1:0] matmul_23_col_select;
  reg [1-1:0] matmul_23_row_select;
  reg [32-1:0] matmul_23_out_col_count;
  reg [32-1:0] matmul_23_out_row_count;
  reg [32-1:0] matmul_23_out_ram_select;
  reg [32-1:0] matmul_23_prev_col_count;
  reg [32-1:0] matmul_23_prev_row_count;
  reg [32-1:0] matmul_23_prev_bat_count;
  reg [32-1:0] matmul_23_prev_och_count;
  reg [1-1:0] matmul_23_prev_row_select;
  reg [32-1:0] matmul_23_stream_act_local_0;
  reg [32-1:0] matmul_23_stream_out_local_val;
  reg [32-1:0] matmul_23_stream_out_local_col;
  wire [32-1:0] matmul_23_stream_out_local;
  assign matmul_23_stream_out_local = matmul_23_stream_out_local_val + matmul_23_stream_out_local_col;
  reg [32-1:0] matmul_23_act_page_comp_offset_0;
  reg [32-1:0] matmul_23_act_page_dma_offset_0;
  reg [32-1:0] matmul_23_filter_page_comp_offset;
  reg [32-1:0] matmul_23_filter_page_dma_offset;
  reg matmul_23_out_page;
  reg [32-1:0] matmul_23_out_page_comp_offset;
  reg [32-1:0] matmul_23_out_page_dma_offset;
  reg [32-1:0] matmul_23_out_laddr_offset;
  reg matmul_23_skip_read_filter;
  reg matmul_23_skip_read_act;
  reg matmul_23_skip_comp;
  reg matmul_23_skip_write_out;
  wire [11-1:0] _dma_read_packed_high_local_size_1306;
  assign _dma_read_packed_high_local_size_1306 = cparam_matmul_23_bias_num >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_1307;
  assign _dma_read_packed_low_local_size_1307 = cparam_matmul_23_bias_num & { 1{ 1'd1 } };
  wire [11-1:0] _dma_read_packed_local_packed_size_1308;
  assign _dma_read_packed_local_packed_size_1308 = (_dma_read_packed_low_local_size_1307 > 0)? _dma_read_packed_high_local_size_1306 + 1 : _dma_read_packed_high_local_size_1306;
  wire [32-1:0] mask_addr_shifted_1309;
  assign mask_addr_shifted_1309 = matmul_23_arg_objaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1310;
  assign mask_addr_masked_1310 = mask_addr_shifted_1309 << 2;
  reg [32-1:0] write_burst_packed_fsm_27;
  localparam write_burst_packed_fsm_27_init = 0;
  reg [10-1:0] write_burst_packed_addr_1311;
  reg [10-1:0] write_burst_packed_stride_1312;
  reg [33-1:0] write_burst_packed_length_1313;
  reg write_burst_packed_done_1314;
  wire [9-1:0] write_burst_packed_ram_addr_1315;
  assign write_burst_packed_ram_addr_1315 = write_burst_packed_addr_1311 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1316;
  assign write_burst_packed_ram_wdata_1316 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l1024_id0_0_1_addr = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1315 : 
                                      ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_210)? write_burst_packed_ram_addr_216 : 'hx;
  assign ram_w16_l1024_id0_0_1_wdata = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1316 : 
                                       ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_210)? write_burst_packed_ram_wdata_217 : 'hx;
  assign ram_w16_l1024_id0_0_1_wenable = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                         ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_210)? 1'd1 : 0;
  assign ram_w16_l1024_id0_0_1_enable = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_210)? 1'd1 : 0;
  wire [9-1:0] write_burst_packed_ram_addr_1317;
  assign write_burst_packed_ram_addr_1317 = write_burst_packed_addr_1311 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1318;
  assign write_burst_packed_ram_wdata_1318 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l1024_id0_1_1_addr = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1317 : 
                                      ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_210)? write_burst_packed_ram_addr_218 : 'hx;
  assign ram_w16_l1024_id0_1_1_wdata = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1318 : 
                                       ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_210)? write_burst_packed_ram_wdata_219 : 'hx;
  assign ram_w16_l1024_id0_1_1_wenable = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                         ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_210)? 1'd1 : 0;
  assign ram_w16_l1024_id0_1_1_enable = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_210)? 1'd1 : 0;
  wire [11-1:0] _dma_read_packed_high_local_size_1319;
  assign _dma_read_packed_high_local_size_1319 = cparam_matmul_23_scale_num >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_1320;
  assign _dma_read_packed_low_local_size_1320 = cparam_matmul_23_scale_num & { 1{ 1'd1 } };
  wire [11-1:0] _dma_read_packed_local_packed_size_1321;
  assign _dma_read_packed_local_packed_size_1321 = (_dma_read_packed_low_local_size_1320 > 0)? _dma_read_packed_high_local_size_1319 + 1 : _dma_read_packed_high_local_size_1319;
  wire [32-1:0] mask_addr_shifted_1322;
  assign mask_addr_shifted_1322 = matmul_23_arg_objaddr_3 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1323;
  assign mask_addr_masked_1323 = mask_addr_shifted_1322 << 2;
  reg [32-1:0] write_burst_packed_fsm_28;
  localparam write_burst_packed_fsm_28_init = 0;
  reg [10-1:0] write_burst_packed_addr_1324;
  reg [10-1:0] write_burst_packed_stride_1325;
  reg [33-1:0] write_burst_packed_length_1326;
  reg write_burst_packed_done_1327;
  wire [9-1:0] write_burst_packed_ram_addr_1328;
  assign write_burst_packed_ram_addr_1328 = write_burst_packed_addr_1324 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1329;
  assign write_burst_packed_ram_wdata_1329 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l1024_id1_0_1_addr = ((write_burst_packed_fsm_28 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1328 : 
                                      ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_220)? write_burst_packed_ram_addr_226 : 'hx;
  assign ram_w16_l1024_id1_0_1_wdata = ((write_burst_packed_fsm_28 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1329 : 
                                       ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_220)? write_burst_packed_ram_wdata_227 : 'hx;
  assign ram_w16_l1024_id1_0_1_wenable = ((write_burst_packed_fsm_28 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                         ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_220)? 1'd1 : 0;
  assign ram_w16_l1024_id1_0_1_enable = ((write_burst_packed_fsm_28 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_220)? 1'd1 : 0;
  wire [9-1:0] write_burst_packed_ram_addr_1330;
  assign write_burst_packed_ram_addr_1330 = write_burst_packed_addr_1324 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1331;
  assign write_burst_packed_ram_wdata_1331 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l1024_id1_1_1_addr = ((write_burst_packed_fsm_28 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1330 : 
                                      ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_220)? write_burst_packed_ram_addr_228 : 'hx;
  assign ram_w16_l1024_id1_1_1_wdata = ((write_burst_packed_fsm_28 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1331 : 
                                       ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_220)? write_burst_packed_ram_wdata_229 : 'hx;
  assign ram_w16_l1024_id1_1_1_wenable = ((write_burst_packed_fsm_28 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                         ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_220)? 1'd1 : 0;
  assign ram_w16_l1024_id1_1_1_enable = ((write_burst_packed_fsm_28 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_220)? 1'd1 : 0;
  wire [14-1:0] _dma_read_packed_high_local_size_1332;
  assign _dma_read_packed_high_local_size_1332 = cparam_matmul_23_filter_read_size >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_1333;
  assign _dma_read_packed_low_local_size_1333 = cparam_matmul_23_filter_read_size & { 1{ 1'd1 } };
  wire [14-1:0] _dma_read_packed_local_packed_size_1334;
  assign _dma_read_packed_local_packed_size_1334 = (_dma_read_packed_low_local_size_1333 > 0)? _dma_read_packed_high_local_size_1332 + 1 : _dma_read_packed_high_local_size_1332;
  wire [32-1:0] mask_addr_shifted_1335;
  assign mask_addr_shifted_1335 = matmul_23_arg_objaddr_1 + matmul_23_filter_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1336;
  assign mask_addr_masked_1336 = mask_addr_shifted_1335 << 2;
  reg [32-1:0] write_burst_packed_fsm_29;
  localparam write_burst_packed_fsm_29_init = 0;
  reg [14-1:0] write_burst_packed_addr_1337;
  reg [14-1:0] write_burst_packed_stride_1338;
  reg [33-1:0] write_burst_packed_length_1339;
  reg write_burst_packed_done_1340;
  wire [13-1:0] write_burst_packed_ram_addr_1341;
  assign write_burst_packed_ram_addr_1341 = write_burst_packed_addr_1337 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1342;
  assign write_burst_packed_ram_wdata_1342 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l16384_id0_0_1_addr = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1341 : 'hx;
  assign ram_w16_l16384_id0_0_1_wdata = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1342 : 'hx;
  assign ram_w16_l16384_id0_0_1_wenable = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l16384_id0_0_1_enable = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [13-1:0] write_burst_packed_ram_addr_1343;
  assign write_burst_packed_ram_addr_1343 = write_burst_packed_addr_1337 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1344;
  assign write_burst_packed_ram_wdata_1344 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l16384_id0_1_1_addr = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1343 : 'hx;
  assign ram_w16_l16384_id0_1_1_wdata = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1344 : 'hx;
  assign ram_w16_l16384_id0_1_1_wenable = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l16384_id0_1_1_enable = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [32-1:0] matmul_23_mux_act_gaddr_0;
  assign matmul_23_mux_act_gaddr_0 = (matmul_23_row_select == 0)? matmul_23_arg_objaddr_0 + (matmul_23_act_base_offset + cparam_matmul_23_act_offset_values_0) : 1'd0;
  wire matmul_23_dma_pad_mask_0;
  assign matmul_23_dma_pad_mask_0 = (matmul_23_row_count + 0 < cparam_matmul_23_pad_row_top) || (matmul_23_row_count + 0 >= cparam_matmul_23_act_num_row + cparam_matmul_23_pad_row_top);
  wire matmul_23_mux_dma_pad_mask_0;
  assign matmul_23_mux_dma_pad_mask_0 = (matmul_23_row_select == 0)? matmul_23_dma_pad_mask_0 : 1'd0;
  wire matmul_23_mux_dma_flag_0;
  assign matmul_23_mux_dma_flag_0 = (matmul_23_prev_row_select == 0)? matmul_23_dma_flag_0 : 1'd0;
  wire [13-1:0] _dma_read_packed_high_local_size_1345;
  assign _dma_read_packed_high_local_size_1345 = cparam_matmul_23_act_read_size >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_1346;
  assign _dma_read_packed_low_local_size_1346 = cparam_matmul_23_act_read_size & { 1{ 1'd1 } };
  wire [13-1:0] _dma_read_packed_local_packed_size_1347;
  assign _dma_read_packed_local_packed_size_1347 = (_dma_read_packed_low_local_size_1346 > 0)? _dma_read_packed_high_local_size_1345 + 1 : _dma_read_packed_high_local_size_1345;
  wire [32-1:0] mask_addr_shifted_1348;
  assign mask_addr_shifted_1348 = matmul_23_mux_act_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1349;
  assign mask_addr_masked_1349 = mask_addr_shifted_1348 << 2;
  reg [32-1:0] write_burst_packed_fsm_30;
  localparam write_burst_packed_fsm_30_init = 0;
  reg [12-1:0] write_burst_packed_addr_1350;
  reg [12-1:0] write_burst_packed_stride_1351;
  reg [33-1:0] write_burst_packed_length_1352;
  reg write_burst_packed_done_1353;
  wire [11-1:0] write_burst_packed_ram_addr_1354;
  assign write_burst_packed_ram_addr_1354 = write_burst_packed_addr_1350 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1355;
  assign write_burst_packed_ram_wdata_1355 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l4096_id0_0_1_addr = ((write_burst_packed_fsm_30 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1354 : 'hx;
  assign ram_w16_l4096_id0_0_1_wdata = ((write_burst_packed_fsm_30 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1355 : 'hx;
  assign ram_w16_l4096_id0_0_1_wenable = ((write_burst_packed_fsm_30 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l4096_id0_0_1_enable = ((write_burst_packed_fsm_30 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [11-1:0] write_burst_packed_ram_addr_1356;
  assign write_burst_packed_ram_addr_1356 = write_burst_packed_addr_1350 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1357;
  assign write_burst_packed_ram_wdata_1357 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l4096_id0_1_1_addr = ((write_burst_packed_fsm_30 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1356 : 'hx;
  assign ram_w16_l4096_id0_1_1_wdata = ((write_burst_packed_fsm_30 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1357 : 'hx;
  assign ram_w16_l4096_id0_1_1_wenable = ((write_burst_packed_fsm_30 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l4096_id0_1_1_enable = ((write_burst_packed_fsm_30 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  reg [32-1:0] matmul_23_comp_fsm;
  localparam matmul_23_comp_fsm_init = 0;
  reg [32-1:0] matmul_23_filter_page_comp_offset_buf;
  reg [32-1:0] matmul_23_act_page_comp_offset_buf_0;
  reg [32-1:0] matmul_23_out_page_comp_offset_buf;
  reg [32-1:0] matmul_23_row_count_buf;
  reg [1-1:0] matmul_23_row_select_buf;
  reg [32-1:0] matmul_23_och_count_buf;
  wire matmul_23_stream_pad_mask_0_0;
  assign matmul_23_stream_pad_mask_0_0 = (matmul_23_col_count + 0 < cparam_matmul_23_pad_col_left) || (matmul_23_col_count + 0 >= cparam_matmul_23_act_num_col + cparam_matmul_23_pad_col_left) || (matmul_23_row_count_buf + 0 < cparam_matmul_23_pad_row_top) || (matmul_23_row_count_buf + 0 >= cparam_matmul_23_act_num_row + cparam_matmul_23_pad_row_top);
  reg [1-1:0] matmul_23_stream_pad_masks;
  wire [13-1:0] stream_matmul_23_parameter_0_data;
  wire [1-1:0] stream_matmul_23_parameter_1_data;
  wire [1-1:0] stream_matmul_23_parameter_2_data;
  wire [1-1:0] stream_matmul_23_parameter_3_data;
  wire [1-1:0] stream_matmul_23_parameter_4_data;
  wire [1-1:0] stream_matmul_23__reduce_reset_data;
  wire [1-1:0] stream_matmul_23_parameter_6_data;
  wire [16-1:0] stream_matmul_23_source_7_data;
  wire [1-1:0] stream_matmul_23_parameter_8_data;
  wire [16-1:0] stream_matmul_23_source_9_data;
  wire [1-1:0] stream_matmul_23_parameter_10_data;
  wire [16-1:0] stream_matmul_23_source_11_data;
  wire [1-1:0] stream_matmul_23_parameter_12_data;
  wire [16-1:0] stream_matmul_23_source_13_data;
  wire [1-1:0] stream_matmul_23_parameter_14_data;
  wire [16-1:0] stream_matmul_23_source_15_data;
  wire [1-1:0] stream_matmul_23_parameter_16_data;
  wire [1-1:0] stream_matmul_23_parameter_17_data;
  wire [1-1:0] stream_matmul_23_parameter_18_data;
  wire [1-1:0] stream_matmul_23_parameter_19_data;
  wire [16-1:0] stream_matmul_23_source_20_data;
  wire [16-1:0] stream_matmul_23_source_21_data;
  reg __stream_matmul_23_stream_ivalid_1;
  reg __stream_matmul_23_stream_ivalid_2;
  reg __stream_matmul_23_stream_ivalid_3;
  reg __stream_matmul_23_stream_ivalid_4;
  reg __stream_matmul_23_stream_ivalid_5;
  reg __stream_matmul_23_stream_ivalid_6;
  reg __stream_matmul_23_stream_ivalid_7;
  reg __stream_matmul_23_stream_ivalid_8;
  reg __stream_matmul_23_stream_ivalid_9;
  reg __stream_matmul_23_stream_ivalid_10;
  reg __stream_matmul_23_stream_ivalid_11;
  reg __stream_matmul_23_stream_ivalid_12;
  reg __stream_matmul_23_stream_ivalid_13;
  reg __stream_matmul_23_stream_ivalid_14;
  reg __stream_matmul_23_stream_ivalid_15;
  reg __stream_matmul_23_stream_ivalid_16;
  reg __stream_matmul_23_stream_ivalid_17;
  reg __stream_matmul_23_stream_ivalid_18;
  reg __stream_matmul_23_stream_ivalid_19;
  reg __stream_matmul_23_stream_ivalid_20;
  reg __stream_matmul_23_stream_ivalid_21;
  reg __stream_matmul_23_stream_ivalid_22;
  reg __stream_matmul_23_stream_ivalid_23;
  reg __stream_matmul_23_stream_ivalid_24;
  reg __stream_matmul_23_stream_ivalid_25;
  reg __stream_matmul_23_stream_ivalid_26;
  reg __stream_matmul_23_stream_ivalid_27;
  reg __stream_matmul_23_stream_ivalid_28;
  reg __stream_matmul_23_stream_ivalid_29;
  wire [16-1:0] _slice_data_975;
  assign _slice_data_975 = stream_matmul_23_source_7_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_976;
  assign _reinterpretcast_src_976 = _slice_data_975;
  wire signed [16-1:0] _reinterpretcast_data_976;
  assign _reinterpretcast_data_976 = _reinterpretcast_src_976;
  wire signed [16-1:0] _cond_data_977;
  assign _cond_data_977 = (stream_matmul_23_parameter_6_data)? _reinterpretcast_data_976 : _reinterpretcast_data_976;
  wire [16-1:0] _slice_data_982;
  assign _slice_data_982 = stream_matmul_23_source_9_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_983;
  assign _reinterpretcast_src_983 = _slice_data_982;
  wire signed [16-1:0] _reinterpretcast_data_983;
  assign _reinterpretcast_data_983 = _reinterpretcast_src_983;
  wire signed [16-1:0] _cond_data_984;
  assign _cond_data_984 = (stream_matmul_23_parameter_8_data)? _reinterpretcast_data_983 : _reinterpretcast_data_983;
  wire [16-1:0] _slice_data_989;
  assign _slice_data_989 = stream_matmul_23_source_11_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_990;
  assign _reinterpretcast_src_990 = _slice_data_989;
  wire [16-1:0] _reinterpretcast_data_990;
  assign _reinterpretcast_data_990 = _reinterpretcast_src_990;
  wire [16-1:0] _cond_data_991;
  assign _cond_data_991 = (stream_matmul_23_parameter_10_data)? _reinterpretcast_data_990 : _reinterpretcast_data_990;
  wire [16-1:0] _slice_data_996;
  assign _slice_data_996 = stream_matmul_23_source_13_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_997;
  assign _reinterpretcast_src_997 = _slice_data_996;
  wire [16-1:0] _reinterpretcast_data_997;
  assign _reinterpretcast_data_997 = _reinterpretcast_src_997;
  wire [16-1:0] _cond_data_998;
  assign _cond_data_998 = (stream_matmul_23_parameter_12_data)? _reinterpretcast_data_997 : _reinterpretcast_data_997;
  wire [16-1:0] _slice_data_1003;
  assign _slice_data_1003 = stream_matmul_23_source_15_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1004;
  assign _reinterpretcast_src_1004 = _slice_data_1003;
  wire [16-1:0] _reinterpretcast_data_1004;
  assign _reinterpretcast_data_1004 = _reinterpretcast_src_1004;
  wire [16-1:0] _cond_data_1005;
  assign _cond_data_1005 = (stream_matmul_23_parameter_14_data)? _reinterpretcast_data_1004 : _reinterpretcast_data_1004;
  reg [1-1:0] _eq_data_1011;
  reg [1-1:0] _eq_data_1015;
  wire [16-1:0] _reinterpretcast_src_1029;
  assign _reinterpretcast_src_1029 = stream_matmul_23_source_21_data;
  wire signed [16-1:0] _reinterpretcast_data_1029;
  assign _reinterpretcast_data_1029 = _reinterpretcast_src_1029;
  wire [1-1:0] _pointer_data_1030;
  assign _pointer_data_1030 = stream_matmul_23_parameter_3_data[1'sd0];
  reg [16-1:0] _plus_data_1035;
  reg [16-1:0] _plus_data_1040;
  reg [16-1:0] _plus_data_1045;
  reg [16-1:0] __delay_data_1401__variable_1010;
  reg [1-1:0] __delay_data_1402_pointer_1030;
  reg signed [16-1:0] __delay_data_1403_reinterpretcast_1029;
  reg [1-1:0] __delay_data_1404__variable_961;
  reg [13-1:0] __delay_data_1425__variable_956;
  reg signed [16-1:0] __delay_data_1436_cond_977;
  reg signed [16-1:0] __delay_data_1453_cond_984;
  wire signed [16-1:0] _cond_data_1013;
  assign _cond_data_1013 = (_eq_data_1011)? __delay_data_1401__variable_1010 : 1'sd0;
  wire signed [16-1:0] _cond_data_1017;
  assign _cond_data_1017 = (_eq_data_1015)? _cond_data_1013 : 1'sd0;
  wire signed [16-1:0] _reinterpretcast_src_1023;
  assign _reinterpretcast_src_1023 = _cond_data_1017;
  wire signed [16-1:0] _reinterpretcast_data_1023;
  assign _reinterpretcast_data_1023 = _reinterpretcast_src_1023;
  wire signed [16-1:0] _cond_data_1033;
  assign _cond_data_1033 = (__delay_data_1402_pointer_1030)? 1'sd0 : _reinterpretcast_data_1023;
  reg [1-1:0] __delay_data_1405__delay_1404__variable_961;
  reg [16-1:0] __delay_data_1415_plus_1040;
  reg [13-1:0] __delay_data_1426__delay_1425__variable_956;
  reg signed [16-1:0] __delay_data_1437__delay_1436_cond_977;
  reg signed [16-1:0] __delay_data_1454__delay_1453_cond_984;
  reg [16-1:0] __delay_data_1471_plus_1045;
  reg [1-1:0] __delay_data_1406__delay_1405__delay_1404__variable_961;
  reg [16-1:0] __delay_data_1416__delay_1415_plus_1040;
  reg [13-1:0] __delay_data_1427__delay_1426__delay_1425__variable_956;
  reg signed [16-1:0] __delay_data_1438__delay_1437__delay_1436_cond_977;
  reg signed [16-1:0] __delay_data_1455__delay_1454__delay_1453_cond_984;
  reg [16-1:0] __delay_data_1472__delay_1471_plus_1045;
  reg [1-1:0] __delay_data_1407__delay_1406__delay_1405____variable_961;
  reg [16-1:0] __delay_data_1417__delay_1416__delay_1415_plus_1040;
  reg [13-1:0] __delay_data_1428__delay_1427__delay_1426____variable_956;
  reg signed [16-1:0] __delay_data_1439__delay_1438__delay_1437__delay_1436_cond_977;
  reg signed [16-1:0] __delay_data_1456__delay_1455__delay_1454__delay_1453_cond_984;
  reg [16-1:0] __delay_data_1473__delay_1472__delay_1471_plus_1045;
  reg [1-1:0] __delay_data_1408__delay_1407__delay_1406____variable_961;
  reg [16-1:0] __delay_data_1418__delay_1417__delay_1416___plus_1040;
  reg [13-1:0] __delay_data_1429__delay_1428__delay_1427____variable_956;
  reg signed [16-1:0] __delay_data_1440__delay_1439__delay_1438__delay_1437___cond_977;
  reg signed [16-1:0] __delay_data_1457__delay_1456__delay_1455__delay_1454___cond_984;
  reg [16-1:0] __delay_data_1474__delay_1473__delay_1472___plus_1045;
  reg [1-1:0] __delay_data_1409__delay_1408__delay_1407____variable_961;
  reg [16-1:0] __delay_data_1419__delay_1418__delay_1417___plus_1040;
  reg [13-1:0] __delay_data_1430__delay_1429__delay_1428____variable_956;
  reg signed [16-1:0] __delay_data_1441__delay_1440__delay_1439__delay_1438___cond_977;
  reg signed [16-1:0] __delay_data_1458__delay_1457__delay_1456__delay_1455___cond_984;
  reg [16-1:0] __delay_data_1475__delay_1474__delay_1473___plus_1045;
  reg [1-1:0] __delay_data_1410__delay_1409__delay_1408____variable_961;
  reg [16-1:0] __delay_data_1420__delay_1419__delay_1418___plus_1040;
  reg [13-1:0] __delay_data_1431__delay_1430__delay_1429____variable_956;
  reg signed [16-1:0] __delay_data_1442__delay_1441__delay_1440__delay_1439___cond_977;
  reg signed [16-1:0] __delay_data_1459__delay_1458__delay_1457__delay_1456___cond_984;
  reg [16-1:0] __delay_data_1476__delay_1475__delay_1474___plus_1045;
  reg [1-1:0] __delay_data_1411__delay_1410__delay_1409____variable_961;
  reg [16-1:0] __delay_data_1421__delay_1420__delay_1419___plus_1040;
  reg [13-1:0] __delay_data_1432__delay_1431__delay_1430____variable_956;
  reg signed [16-1:0] __delay_data_1443__delay_1442__delay_1441__delay_1440___cond_977;
  reg signed [16-1:0] __delay_data_1460__delay_1459__delay_1458__delay_1457___cond_984;
  reg [16-1:0] __delay_data_1477__delay_1476__delay_1475___plus_1045;
  reg [1-1:0] __delay_data_1412__delay_1411__delay_1410____variable_961;
  reg [16-1:0] __delay_data_1422__delay_1421__delay_1420___plus_1040;
  reg [13-1:0] __delay_data_1433__delay_1432__delay_1431____variable_956;
  reg signed [16-1:0] __delay_data_1444__delay_1443__delay_1442__delay_1441___cond_977;
  reg signed [16-1:0] __delay_data_1461__delay_1460__delay_1459__delay_1458___cond_984;
  reg [16-1:0] __delay_data_1478__delay_1477__delay_1476___plus_1045;
  reg [1-1:0] __delay_data_1413__delay_1412__delay_1411____variable_961;
  reg [16-1:0] __delay_data_1423__delay_1422__delay_1421___plus_1040;
  reg [13-1:0] __delay_data_1434__delay_1433__delay_1432____variable_956;
  reg signed [16-1:0] __delay_data_1445__delay_1444__delay_1443__delay_1442___cond_977;
  reg signed [16-1:0] __delay_data_1462__delay_1461__delay_1460__delay_1459___cond_984;
  reg [16-1:0] __delay_data_1479__delay_1478__delay_1477___plus_1045;
  wire signed [32-1:0] __substreamoutput_data_1036;
  assign __substreamoutput_data_1036 = mul_8_z_data;
  reg signed [64-1:0] __variable_wdata_44;
  assign add_tree_2_var0_data = __variable_wdata_44;
  assign _add_tree_2_is_root = ((_stream_matmul_23_busy)? 0 : 1) && 1;
  assign _add_tree_2_stream_oready = ((_stream_matmul_23_busy)? _stream_matmul_23_stream_oready : 1) && _add_tree_2_stream_internal_oready;
  reg [1-1:0] __delay_data_1414__delay_1413__delay_1412____variable_961;
  reg [16-1:0] __delay_data_1424__delay_1423__delay_1422___plus_1040;
  reg [13-1:0] __delay_data_1435__delay_1434__delay_1433____variable_956;
  reg signed [16-1:0] __delay_data_1446__delay_1445__delay_1444__delay_1443___cond_977;
  reg signed [16-1:0] __delay_data_1463__delay_1462__delay_1461__delay_1460___cond_984;
  reg [16-1:0] __delay_data_1480__delay_1479__delay_1478___plus_1045;
  wire signed [64-1:0] __substreamoutput_data_1038;
  assign __substreamoutput_data_1038 = add_tree_2_sum_data;
  reg signed [16-1:0] __delay_data_1447__delay_1446__delay_1445__delay_1444___cond_977;
  reg signed [16-1:0] __delay_data_1464__delay_1463__delay_1462__delay_1461___cond_984;
  reg [16-1:0] __delay_data_1481__delay_1480__delay_1479___plus_1045;
  reg signed [16-1:0] __delay_data_1448__delay_1447__delay_1446__delay_1445___cond_977;
  reg signed [16-1:0] __delay_data_1465__delay_1464__delay_1463__delay_1462___cond_984;
  reg [16-1:0] __delay_data_1482__delay_1481__delay_1480___plus_1045;
  reg signed [16-1:0] __delay_data_1449__delay_1448__delay_1447__delay_1446___cond_977;
  reg signed [16-1:0] __delay_data_1466__delay_1465__delay_1464__delay_1463___cond_984;
  reg [16-1:0] __delay_data_1483__delay_1482__delay_1481___plus_1045;
  reg signed [16-1:0] __delay_data_1450__delay_1449__delay_1448__delay_1447___cond_977;
  reg signed [16-1:0] __delay_data_1467__delay_1466__delay_1465__delay_1464___cond_984;
  reg [16-1:0] __delay_data_1484__delay_1483__delay_1482___plus_1045;
  reg signed [16-1:0] __delay_data_1451__delay_1450__delay_1449__delay_1448___cond_977;
  reg signed [16-1:0] __delay_data_1468__delay_1467__delay_1466__delay_1465___cond_984;
  reg [16-1:0] __delay_data_1485__delay_1484__delay_1483___plus_1045;
  reg signed [16-1:0] __delay_data_1452__delay_1451__delay_1450__delay_1449___cond_977;
  reg signed [16-1:0] __delay_data_1469__delay_1468__delay_1467__delay_1466___cond_984;
  reg [16-1:0] __delay_data_1486__delay_1485__delay_1484___plus_1045;
  wire signed [64-1:0] __substreamoutput_data_1041;
  assign __substreamoutput_data_1041 = acc_0_sum_data;
  wire [1-1:0] __substreamoutput_data_1042;
  assign __substreamoutput_data_1042 = acc_0_valid_data;
  reg signed [64-1:0] _plus_data_1043;
  reg signed [16-1:0] __delay_data_1470__delay_1469__delay_1468__delay_1467___cond_984;
  reg [16-1:0] __delay_data_1487__delay_1486__delay_1485___plus_1045;
  reg [1-1:0] __delay_data_1489__substreamoutput_1042;
  assign _stream_matmul_23_stream_internal_oready = ((_stream_matmul_23_busy)? _mul_rshift_round_clip_6_stream_internal_oready : 1) && (((_stream_matmul_23_busy)? _acc_0_stream_internal_oready : 1) && (((_stream_matmul_23_busy)? _add_tree_2_stream_internal_oready : 1) && (((_stream_matmul_23_busy)? _mul_8_stream_internal_oready : 1) && 1)));
  reg [1-1:0] __delay_data_1490__delay_1489__substreamoutput_1042;
  reg [1-1:0] __delay_data_1491__delay_1490____substreamoutput_1042;
  reg [1-1:0] __delay_data_1492__delay_1491____substreamoutput_1042;
  reg [1-1:0] __delay_data_1493__delay_1492____substreamoutput_1042;
  reg [1-1:0] __delay_data_1494__delay_1493____substreamoutput_1042;
  reg [1-1:0] __delay_data_1495__delay_1494____substreamoutput_1042;
  reg [1-1:0] __delay_data_1496__delay_1495____substreamoutput_1042;
  reg [1-1:0] __delay_data_1497__delay_1496____substreamoutput_1042;
  reg [1-1:0] __delay_data_1498__delay_1497____substreamoutput_1042;
  wire signed [16-1:0] __substreamoutput_data_1046;
  assign __substreamoutput_data_1046 = mul_rshift_round_clip_6_z_data;
  reg [1-1:0] _greaterthan_data_1048;
  reg signed [16-1:0] __delay_data_1488__substreamoutput_1046;
  reg [1-1:0] __delay_data_1499__delay_1498____substreamoutput_1042;
  reg signed [16-1:0] _cond_data_1050;
  reg [1-1:0] __delay_data_1500__delay_1499____substreamoutput_1042;
  wire signed [16-1:0] _reinterpretcast_src_1051;
  assign _reinterpretcast_src_1051 = _cond_data_1050;
  wire signed [16-1:0] _reinterpretcast_data_1051;
  assign _reinterpretcast_data_1051 = _reinterpretcast_src_1051;
  wire signed [16-1:0] stream_matmul_23_sink_26_data;
  assign stream_matmul_23_sink_26_data = _reinterpretcast_data_1051;
  wire [1-1:0] stream_matmul_23_sink_27_data;
  assign stream_matmul_23_sink_27_data = __delay_data_1500__delay_1499____substreamoutput_1042;
  wire _set_flag_1358;
  assign _set_flag_1358 = matmul_23_comp_fsm == 3;
  reg [13-1:0] __variable_wdata_956;
  assign stream_matmul_23_parameter_0_data = __variable_wdata_956;
  wire _set_flag_1359;
  assign _set_flag_1359 = matmul_23_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_957;
  assign stream_matmul_23_parameter_1_data = __variable_wdata_957;
  wire _set_flag_1360;
  assign _set_flag_1360 = matmul_23_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_958;
  assign stream_matmul_23_parameter_2_data = __variable_wdata_958;
  wire _set_flag_1361;
  assign _set_flag_1361 = matmul_23_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_959;
  assign stream_matmul_23_parameter_3_data = __variable_wdata_959;
  wire _set_flag_1362;
  assign _set_flag_1362 = matmul_23_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_960;
  assign stream_matmul_23_parameter_4_data = __variable_wdata_960;
  wire _set_flag_1363;
  assign _set_flag_1363 = matmul_23_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_971;
  assign stream_matmul_23_parameter_6_data = __variable_wdata_971;
  reg [32-1:0] _source_stream_matmul_23_source_7_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_23_source_7_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_23_source_7_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_23_source_7_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_23_source_7_pat_size_0;
  reg [33-1:0] _source_stream_matmul_23_source_7_pat_size_1;
  reg [33-1:0] _source_stream_matmul_23_source_7_pat_size_2;
  reg [33-1:0] _source_stream_matmul_23_source_7_pat_size_3;
  reg [32-1:0] _source_stream_matmul_23_source_7_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_23_source_7_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_23_source_7_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_23_source_7_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_23_source_7_pat_count_0;
  reg [33-1:0] _source_stream_matmul_23_source_7_pat_count_1;
  reg [33-1:0] _source_stream_matmul_23_source_7_pat_count_2;
  reg [33-1:0] _source_stream_matmul_23_source_7_pat_count_3;
  reg [33-1:0] _source_stream_matmul_23_source_7_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_23_source_7_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_23_source_7_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_23_source_7_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_23_source_7_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_23_source_7_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_23_source_7_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_23_source_7_pat_stride_buf_3;
  wire _set_flag_1364;
  assign _set_flag_1364 = matmul_23_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_1365;
  assign read_rtl_bank_1365 = _stream_matmul_23_source_7_source_ram_raddr;
  reg [1-1:0] _tmp_1366;
  assign ram_w16_l1024_id0_0_0_addr = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_7_source_ram_renable && (_stream_matmul_23_source_7_source_sel == 1))? _stream_matmul_23_source_7_source_ram_raddr >> 1 : 
                                      (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3))? _stream_conv2d_4_source_20_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id0_0_0_enable = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_7_source_ram_renable && (_stream_matmul_23_source_7_source_sel == 1))? 1'd1 : 
                                        (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1367 = 1;
  wire [_tmp_1367-1:0] _tmp_1368;
  assign _tmp_1368 = _stream_matmul_23_stream_oready && _stream_matmul_23_source_7_source_ram_renable && (_stream_matmul_23_source_7_source_sel == 1);
  reg [_tmp_1367-1:0] __tmp_1368_1;
  assign ram_w16_l1024_id0_1_0_addr = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_7_source_ram_renable && (_stream_matmul_23_source_7_source_sel == 1))? _stream_matmul_23_source_7_source_ram_raddr >> 1 : 
                                      (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3))? _stream_conv2d_4_source_20_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id0_1_0_enable = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_7_source_ram_renable && (_stream_matmul_23_source_7_source_sel == 1))? 1'd1 : 
                                        (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1369 = 1;
  wire [_tmp_1369-1:0] _tmp_1370;
  assign _tmp_1370 = _stream_matmul_23_stream_oready && _stream_matmul_23_source_7_source_ram_renable && (_stream_matmul_23_source_7_source_sel == 1);
  reg [_tmp_1369-1:0] __tmp_1370_1;
  wire signed [16-1:0] read_rtl_rdata_1371;
  wire read_rtl_rvalid_1372;
  assign read_rtl_rdata_1371 = (_tmp_1366 == 0)? ram_w16_l1024_id0_0_0_rdata : 
                               (_tmp_1366 == 1)? ram_w16_l1024_id0_1_0_rdata : 0;
  assign read_rtl_rvalid_1372 = __tmp_1368_1;
  assign _stream_matmul_23_source_7_source_ram_rdata = (_stream_matmul_23_source_7_source_sel == 1)? read_rtl_rdata_1371 : 'hx;
  reg [16-1:0] __variable_wdata_972;
  assign stream_matmul_23_source_7_data = __variable_wdata_972;
  reg [32-1:0] _stream_matmul_23_source_7_source_pat_fsm_0;
  localparam _stream_matmul_23_source_7_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_matmul_23_source_7_source_pat_all_offset;
  assign _stream_matmul_23_source_7_source_pat_all_offset = _stream_matmul_23_source_7_source_offset_buf + _source_stream_matmul_23_source_7_pat_cur_offset_0 + _source_stream_matmul_23_source_7_pat_cur_offset_1 + _source_stream_matmul_23_source_7_pat_cur_offset_2 + _source_stream_matmul_23_source_7_pat_cur_offset_3;
  wire _set_flag_1373;
  assign _set_flag_1373 = matmul_23_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_978;
  assign stream_matmul_23_parameter_8_data = __variable_wdata_978;
  reg [32-1:0] _source_stream_matmul_23_source_9_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_23_source_9_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_23_source_9_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_23_source_9_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_23_source_9_pat_size_0;
  reg [33-1:0] _source_stream_matmul_23_source_9_pat_size_1;
  reg [33-1:0] _source_stream_matmul_23_source_9_pat_size_2;
  reg [33-1:0] _source_stream_matmul_23_source_9_pat_size_3;
  reg [32-1:0] _source_stream_matmul_23_source_9_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_23_source_9_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_23_source_9_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_23_source_9_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_23_source_9_pat_count_0;
  reg [33-1:0] _source_stream_matmul_23_source_9_pat_count_1;
  reg [33-1:0] _source_stream_matmul_23_source_9_pat_count_2;
  reg [33-1:0] _source_stream_matmul_23_source_9_pat_count_3;
  reg [33-1:0] _source_stream_matmul_23_source_9_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_23_source_9_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_23_source_9_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_23_source_9_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_23_source_9_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_23_source_9_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_23_source_9_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_23_source_9_pat_stride_buf_3;
  wire _set_flag_1374;
  assign _set_flag_1374 = matmul_23_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_1375;
  assign read_rtl_bank_1375 = _stream_matmul_23_source_9_source_ram_raddr;
  reg [1-1:0] _tmp_1376;
  assign ram_w16_l1024_id1_0_0_addr = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_9_source_ram_renable && (_stream_matmul_23_source_9_source_sel == 2))? _stream_matmul_23_source_9_source_ram_raddr >> 1 : 
                                      (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4))? _stream_conv2d_4_source_21_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id1_0_0_enable = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_9_source_ram_renable && (_stream_matmul_23_source_9_source_sel == 2))? 1'd1 : 
                                        (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4))? 1'd1 : 0;
  localparam _tmp_1377 = 1;
  wire [_tmp_1377-1:0] _tmp_1378;
  assign _tmp_1378 = _stream_matmul_23_stream_oready && _stream_matmul_23_source_9_source_ram_renable && (_stream_matmul_23_source_9_source_sel == 2);
  reg [_tmp_1377-1:0] __tmp_1378_1;
  assign ram_w16_l1024_id1_1_0_addr = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_9_source_ram_renable && (_stream_matmul_23_source_9_source_sel == 2))? _stream_matmul_23_source_9_source_ram_raddr >> 1 : 
                                      (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4))? _stream_conv2d_4_source_21_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l1024_id1_1_0_enable = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_9_source_ram_renable && (_stream_matmul_23_source_9_source_sel == 2))? 1'd1 : 
                                        (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4))? 1'd1 : 0;
  localparam _tmp_1379 = 1;
  wire [_tmp_1379-1:0] _tmp_1380;
  assign _tmp_1380 = _stream_matmul_23_stream_oready && _stream_matmul_23_source_9_source_ram_renable && (_stream_matmul_23_source_9_source_sel == 2);
  reg [_tmp_1379-1:0] __tmp_1380_1;
  wire signed [16-1:0] read_rtl_rdata_1381;
  wire read_rtl_rvalid_1382;
  assign read_rtl_rdata_1381 = (_tmp_1376 == 0)? ram_w16_l1024_id1_0_0_rdata : 
                               (_tmp_1376 == 1)? ram_w16_l1024_id1_1_0_rdata : 0;
  assign read_rtl_rvalid_1382 = __tmp_1378_1;
  assign _stream_matmul_23_source_9_source_ram_rdata = (_stream_matmul_23_source_9_source_sel == 2)? read_rtl_rdata_1381 : 'hx;
  reg [16-1:0] __variable_wdata_979;
  assign stream_matmul_23_source_9_data = __variable_wdata_979;
  reg [32-1:0] _stream_matmul_23_source_9_source_pat_fsm_1;
  localparam _stream_matmul_23_source_9_source_pat_fsm_1_init = 0;
  wire [32-1:0] _stream_matmul_23_source_9_source_pat_all_offset;
  assign _stream_matmul_23_source_9_source_pat_all_offset = _stream_matmul_23_source_9_source_offset_buf + _source_stream_matmul_23_source_9_pat_cur_offset_0 + _source_stream_matmul_23_source_9_pat_cur_offset_1 + _source_stream_matmul_23_source_9_pat_cur_offset_2 + _source_stream_matmul_23_source_9_pat_cur_offset_3;
  wire _set_flag_1383;
  assign _set_flag_1383 = matmul_23_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_985;
  assign stream_matmul_23_parameter_10_data = __variable_wdata_985;
  wire _set_flag_1384;
  assign _set_flag_1384 = matmul_23_comp_fsm == 3;
  reg [16-1:0] __variable_wdata_986;
  assign stream_matmul_23_source_11_data = __variable_wdata_986;
  wire _set_flag_1385;
  assign _set_flag_1385 = matmul_23_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_992;
  assign stream_matmul_23_parameter_12_data = __variable_wdata_992;
  wire _set_flag_1386;
  assign _set_flag_1386 = matmul_23_comp_fsm == 3;
  reg [16-1:0] __variable_wdata_993;
  assign stream_matmul_23_source_13_data = __variable_wdata_993;
  wire _set_flag_1387;
  assign _set_flag_1387 = matmul_23_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_999;
  assign stream_matmul_23_parameter_14_data = __variable_wdata_999;
  wire _set_flag_1388;
  assign _set_flag_1388 = matmul_23_comp_fsm == 3;
  reg [16-1:0] __variable_wdata_1000;
  assign stream_matmul_23_source_15_data = __variable_wdata_1000;
  wire _set_flag_1389;
  assign _set_flag_1389 = matmul_23_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1006;
  assign stream_matmul_23_parameter_16_data = __variable_wdata_1006;
  wire _set_flag_1390;
  assign _set_flag_1390 = matmul_23_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1007;
  assign stream_matmul_23_parameter_17_data = __variable_wdata_1007;
  wire _set_flag_1391;
  assign _set_flag_1391 = matmul_23_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1008;
  assign stream_matmul_23_parameter_18_data = __variable_wdata_1008;
  wire _set_flag_1392;
  assign _set_flag_1392 = matmul_23_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1009;
  assign stream_matmul_23_parameter_19_data = __variable_wdata_1009;
  reg [32-1:0] _source_stream_matmul_23_source_20_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_23_source_20_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_23_source_20_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_23_source_20_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_23_source_20_pat_size_0;
  reg [33-1:0] _source_stream_matmul_23_source_20_pat_size_1;
  reg [33-1:0] _source_stream_matmul_23_source_20_pat_size_2;
  reg [33-1:0] _source_stream_matmul_23_source_20_pat_size_3;
  reg [32-1:0] _source_stream_matmul_23_source_20_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_23_source_20_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_23_source_20_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_23_source_20_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_23_source_20_pat_count_0;
  reg [33-1:0] _source_stream_matmul_23_source_20_pat_count_1;
  reg [33-1:0] _source_stream_matmul_23_source_20_pat_count_2;
  reg [33-1:0] _source_stream_matmul_23_source_20_pat_count_3;
  reg [33-1:0] _source_stream_matmul_23_source_20_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_23_source_20_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_23_source_20_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_23_source_20_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_23_source_20_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_23_source_20_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_23_source_20_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_23_source_20_pat_stride_buf_3;
  wire _set_flag_1393;
  assign _set_flag_1393 = matmul_23_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_1394;
  assign read_rtl_bank_1394 = _stream_matmul_23_source_20_source_ram_raddr;
  reg [1-1:0] _tmp_1395;
  assign ram_w16_l4096_id0_0_0_addr = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_20_source_ram_renable && (_stream_matmul_23_source_20_source_sel == 3))? _stream_matmul_23_source_20_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l4096_id0_0_0_enable = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_20_source_ram_renable && (_stream_matmul_23_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1396 = 1;
  wire [_tmp_1396-1:0] _tmp_1397;
  assign _tmp_1397 = _stream_matmul_23_stream_oready && _stream_matmul_23_source_20_source_ram_renable && (_stream_matmul_23_source_20_source_sel == 3);
  reg [_tmp_1396-1:0] __tmp_1397_1;
  assign ram_w16_l4096_id0_1_0_addr = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_20_source_ram_renable && (_stream_matmul_23_source_20_source_sel == 3))? _stream_matmul_23_source_20_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l4096_id0_1_0_enable = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_20_source_ram_renable && (_stream_matmul_23_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1398 = 1;
  wire [_tmp_1398-1:0] _tmp_1399;
  assign _tmp_1399 = _stream_matmul_23_stream_oready && _stream_matmul_23_source_20_source_ram_renable && (_stream_matmul_23_source_20_source_sel == 3);
  reg [_tmp_1398-1:0] __tmp_1399_1;
  wire signed [16-1:0] read_rtl_rdata_1400;
  wire read_rtl_rvalid_1401;
  assign read_rtl_rdata_1400 = (_tmp_1395 == 0)? ram_w16_l4096_id0_0_0_rdata : 
                               (_tmp_1395 == 1)? ram_w16_l4096_id0_1_0_rdata : 0;
  assign read_rtl_rvalid_1401 = __tmp_1397_1;
  assign _stream_matmul_23_source_20_source_ram_rdata = (_stream_matmul_23_source_20_source_sel == 3)? read_rtl_rdata_1400 : 'hx;
  reg [16-1:0] __variable_wdata_1010;
  assign stream_matmul_23_source_20_data = __variable_wdata_1010;
  reg [32-1:0] _stream_matmul_23_source_20_source_pat_fsm_2;
  localparam _stream_matmul_23_source_20_source_pat_fsm_2_init = 0;
  wire [32-1:0] _stream_matmul_23_source_20_source_pat_all_offset;
  assign _stream_matmul_23_source_20_source_pat_all_offset = _stream_matmul_23_source_20_source_offset_buf + _source_stream_matmul_23_source_20_pat_cur_offset_0 + _source_stream_matmul_23_source_20_pat_cur_offset_1 + _source_stream_matmul_23_source_20_pat_cur_offset_2 + _source_stream_matmul_23_source_20_pat_cur_offset_3;
  reg [32-1:0] _source_stream_matmul_23_source_21_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_23_source_21_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_23_source_21_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_23_source_21_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_23_source_21_pat_size_0;
  reg [33-1:0] _source_stream_matmul_23_source_21_pat_size_1;
  reg [33-1:0] _source_stream_matmul_23_source_21_pat_size_2;
  reg [33-1:0] _source_stream_matmul_23_source_21_pat_size_3;
  reg [32-1:0] _source_stream_matmul_23_source_21_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_23_source_21_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_23_source_21_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_23_source_21_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_23_source_21_pat_count_0;
  reg [33-1:0] _source_stream_matmul_23_source_21_pat_count_1;
  reg [33-1:0] _source_stream_matmul_23_source_21_pat_count_2;
  reg [33-1:0] _source_stream_matmul_23_source_21_pat_count_3;
  reg [33-1:0] _source_stream_matmul_23_source_21_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_23_source_21_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_23_source_21_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_23_source_21_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_23_source_21_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_23_source_21_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_23_source_21_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_23_source_21_pat_stride_buf_3;
  wire _set_flag_1402;
  assign _set_flag_1402 = matmul_23_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_1403;
  assign read_rtl_bank_1403 = _stream_matmul_23_source_21_source_ram_raddr;
  reg [1-1:0] _tmp_1404;
  assign ram_w16_l16384_id0_0_0_addr = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_21_source_ram_renable && (_stream_matmul_23_source_21_source_sel == 4))? _stream_matmul_23_source_21_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l16384_id0_0_0_enable = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_21_source_ram_renable && (_stream_matmul_23_source_21_source_sel == 4))? 1'd1 : 0;
  localparam _tmp_1405 = 1;
  wire [_tmp_1405-1:0] _tmp_1406;
  assign _tmp_1406 = _stream_matmul_23_stream_oready && _stream_matmul_23_source_21_source_ram_renable && (_stream_matmul_23_source_21_source_sel == 4);
  reg [_tmp_1405-1:0] __tmp_1406_1;
  assign ram_w16_l16384_id0_1_0_addr = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_21_source_ram_renable && (_stream_matmul_23_source_21_source_sel == 4))? _stream_matmul_23_source_21_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l16384_id0_1_0_enable = (_stream_matmul_23_stream_oready && _stream_matmul_23_source_21_source_ram_renable && (_stream_matmul_23_source_21_source_sel == 4))? 1'd1 : 0;
  localparam _tmp_1407 = 1;
  wire [_tmp_1407-1:0] _tmp_1408;
  assign _tmp_1408 = _stream_matmul_23_stream_oready && _stream_matmul_23_source_21_source_ram_renable && (_stream_matmul_23_source_21_source_sel == 4);
  reg [_tmp_1407-1:0] __tmp_1408_1;
  wire signed [16-1:0] read_rtl_rdata_1409;
  wire read_rtl_rvalid_1410;
  assign read_rtl_rdata_1409 = (_tmp_1404 == 0)? ram_w16_l16384_id0_0_0_rdata : 
                               (_tmp_1404 == 1)? ram_w16_l16384_id0_1_0_rdata : 0;
  assign read_rtl_rvalid_1410 = __tmp_1406_1;
  assign _stream_matmul_23_source_21_source_ram_rdata = (_stream_matmul_23_source_21_source_sel == 4)? read_rtl_rdata_1409 : 'hx;
  reg [16-1:0] __variable_wdata_1024;
  assign stream_matmul_23_source_21_data = __variable_wdata_1024;
  reg [32-1:0] _stream_matmul_23_source_21_source_pat_fsm_3;
  localparam _stream_matmul_23_source_21_source_pat_fsm_3_init = 0;
  wire [32-1:0] _stream_matmul_23_source_21_source_pat_all_offset;
  assign _stream_matmul_23_source_21_source_pat_all_offset = _stream_matmul_23_source_21_source_offset_buf + _source_stream_matmul_23_source_21_pat_cur_offset_0 + _source_stream_matmul_23_source_21_pat_cur_offset_1 + _source_stream_matmul_23_source_21_pat_cur_offset_2 + _source_stream_matmul_23_source_21_pat_cur_offset_3;
  wire _set_flag_1411;
  assign _set_flag_1411 = matmul_23_comp_fsm == 3;
  reg _tmp_1412;
  reg _tmp_1413;
  reg _tmp_1414;
  reg _tmp_1415;
  reg _tmp_1416;
  reg _tmp_1417;
  reg _tmp_1418;
  reg _tmp_1419;
  reg _tmp_1420;
  reg _tmp_1421;
  reg _tmp_1422;
  reg _tmp_1423;
  reg _tmp_1424;
  reg _tmp_1425;
  reg _tmp_1426;
  reg _tmp_1427;
  reg _tmp_1428;
  reg _tmp_1429;
  reg _tmp_1430;
  reg _tmp_1431;
  reg _tmp_1432;
  reg _tmp_1433;
  reg _tmp_1434;
  reg _tmp_1435;
  reg _tmp_1436;
  reg _tmp_1437;
  reg _tmp_1438;
  reg _tmp_1439;
  reg _tmp_1440;
  reg _tmp_1441;
  reg _tmp_1442;
  localparam _tmp_1443 = 33;
  wire [_tmp_1443-1:0] _tmp_1444;
  assign _tmp_1444 = matmul_23_stream_out_local + matmul_23_out_page_comp_offset_buf;
  reg [_tmp_1443-1:0] _tmp_1445;
  reg [_tmp_1443-1:0] _tmp_1446;
  reg [_tmp_1443-1:0] _tmp_1447;
  reg [_tmp_1443-1:0] _tmp_1448;
  reg [_tmp_1443-1:0] _tmp_1449;
  reg [_tmp_1443-1:0] _tmp_1450;
  reg [_tmp_1443-1:0] _tmp_1451;
  reg [_tmp_1443-1:0] _tmp_1452;
  reg [_tmp_1443-1:0] _tmp_1453;
  reg [_tmp_1443-1:0] _tmp_1454;
  reg [_tmp_1443-1:0] _tmp_1455;
  reg [_tmp_1443-1:0] _tmp_1456;
  reg [_tmp_1443-1:0] _tmp_1457;
  reg [_tmp_1443-1:0] _tmp_1458;
  reg [_tmp_1443-1:0] _tmp_1459;
  reg [_tmp_1443-1:0] _tmp_1460;
  reg [_tmp_1443-1:0] _tmp_1461;
  reg [_tmp_1443-1:0] _tmp_1462;
  reg [_tmp_1443-1:0] _tmp_1463;
  reg [_tmp_1443-1:0] _tmp_1464;
  reg [_tmp_1443-1:0] _tmp_1465;
  reg [_tmp_1443-1:0] _tmp_1466;
  reg [_tmp_1443-1:0] _tmp_1467;
  reg [_tmp_1443-1:0] _tmp_1468;
  reg [_tmp_1443-1:0] _tmp_1469;
  reg [_tmp_1443-1:0] _tmp_1470;
  reg [_tmp_1443-1:0] _tmp_1471;
  reg [_tmp_1443-1:0] _tmp_1472;
  reg [_tmp_1443-1:0] _tmp_1473;
  reg [_tmp_1443-1:0] _tmp_1474;
  reg [_tmp_1443-1:0] _tmp_1475;
  reg [32-1:0] _tmp_1476;
  reg [32-1:0] _tmp_1477;
  reg [32-1:0] _tmp_1478;
  reg [32-1:0] _tmp_1479;
  reg [32-1:0] _tmp_1480;
  reg [32-1:0] _tmp_1481;
  reg [32-1:0] _tmp_1482;
  reg [32-1:0] _tmp_1483;
  reg [32-1:0] _tmp_1484;
  reg [32-1:0] _tmp_1485;
  reg [32-1:0] _tmp_1486;
  reg [32-1:0] _tmp_1487;
  reg [32-1:0] _tmp_1488;
  reg [32-1:0] _tmp_1489;
  reg [32-1:0] _tmp_1490;
  reg [32-1:0] _tmp_1491;
  reg [32-1:0] _tmp_1492;
  reg [32-1:0] _tmp_1493;
  reg [32-1:0] _tmp_1494;
  reg [32-1:0] _tmp_1495;
  reg [32-1:0] _tmp_1496;
  reg [32-1:0] _tmp_1497;
  reg [32-1:0] _tmp_1498;
  reg [32-1:0] _tmp_1499;
  reg [32-1:0] _tmp_1500;
  reg [32-1:0] _tmp_1501;
  reg [32-1:0] _tmp_1502;
  reg [32-1:0] _tmp_1503;
  reg [32-1:0] _tmp_1504;
  reg [32-1:0] _tmp_1505;
  reg [32-1:0] _tmp_1506;
  wire [1-1:0] write_rtl_bank_1507;
  assign write_rtl_bank_1507 = _stream_matmul_23_sink_26_sink_waddr;
  assign ram_w16_l512_id0_0_0_addr = (_stream_matmul_23_stream_oready && _stream_matmul_23_sink_26_sink_wenable && (_stream_matmul_23_sink_26_sink_sel == 5) && (write_rtl_bank_1507 == 0))? _stream_matmul_23_sink_26_sink_waddr >> 1 : 
                                     (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 0))? _stream_conv2d_4_sink_50_sink_waddr >> 1 : 'hx;
  assign ram_w16_l512_id0_0_0_wdata = (_stream_matmul_23_stream_oready && _stream_matmul_23_sink_26_sink_wenable && (_stream_matmul_23_sink_26_sink_sel == 5) && (write_rtl_bank_1507 == 0))? _stream_matmul_23_sink_26_sink_wdata : 
                                      (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 0))? _stream_conv2d_4_sink_50_sink_wdata : 'hx;
  assign ram_w16_l512_id0_0_0_wenable = (_stream_matmul_23_stream_oready && _stream_matmul_23_sink_26_sink_wenable && (_stream_matmul_23_sink_26_sink_sel == 5) && (write_rtl_bank_1507 == 0))? 1'd1 : 
                                        (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 0))? 1'd1 : 0;
  assign ram_w16_l512_id0_0_0_enable = (_stream_matmul_23_stream_oready && _stream_matmul_23_sink_26_sink_wenable && (_stream_matmul_23_sink_26_sink_sel == 5) && (write_rtl_bank_1507 == 0))? 1'd1 : 
                                       (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 0))? 1'd1 : 0;
  assign ram_w16_l512_id0_1_0_addr = (_stream_matmul_23_stream_oready && _stream_matmul_23_sink_26_sink_wenable && (_stream_matmul_23_sink_26_sink_sel == 5) && (write_rtl_bank_1507 == 1))? _stream_matmul_23_sink_26_sink_waddr >> 1 : 
                                     (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 1))? _stream_conv2d_4_sink_50_sink_waddr >> 1 : 'hx;
  assign ram_w16_l512_id0_1_0_wdata = (_stream_matmul_23_stream_oready && _stream_matmul_23_sink_26_sink_wenable && (_stream_matmul_23_sink_26_sink_sel == 5) && (write_rtl_bank_1507 == 1))? _stream_matmul_23_sink_26_sink_wdata : 
                                      (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 1))? _stream_conv2d_4_sink_50_sink_wdata : 'hx;
  assign ram_w16_l512_id0_1_0_wenable = (_stream_matmul_23_stream_oready && _stream_matmul_23_sink_26_sink_wenable && (_stream_matmul_23_sink_26_sink_sel == 5) && (write_rtl_bank_1507 == 1))? 1'd1 : 
                                        (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 1))? 1'd1 : 0;
  assign ram_w16_l512_id0_1_0_enable = (_stream_matmul_23_stream_oready && _stream_matmul_23_sink_26_sink_wenable && (_stream_matmul_23_sink_26_sink_sel == 5) && (write_rtl_bank_1507 == 1))? 1'd1 : 
                                       (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 1))? 1'd1 : 0;
  reg [32-1:0] _stream_matmul_23_sink_26_sink_fsm_4;
  localparam _stream_matmul_23_sink_26_sink_fsm_4_init = 0;
  wire _set_flag_1508;
  assign _set_flag_1508 = matmul_23_comp_fsm == 4;
  assign _stream_matmul_23_run_flag = (_set_flag_1508)? 1 : 0;
  reg _tmp_1509;
  reg _tmp_1510;
  reg _tmp_1511;
  assign _add_tree_2_source_stop = _add_tree_2_stream_oready && 1'd0;
  reg _tmp_1512;
  reg _tmp_1513;
  assign _add_tree_2_sink_start = _tmp_1513;
  reg _tmp_1514;
  reg _tmp_1515;
  assign _add_tree_2_sink_stop = _tmp_1515;
  reg _tmp_1516;
  reg _tmp_1517;
  assign _add_tree_2_sink_busy = _tmp_1517;
  reg _tmp_1518;
  assign _add_tree_2_busy = _add_tree_2_source_busy || _add_tree_2_sink_busy || _add_tree_2_busy_reg;
  reg _tmp_1519;
  reg _tmp_1520;
  reg _tmp_1521;
  reg _tmp_1522;
  reg _tmp_1523;
  reg _tmp_1524;
  reg [1-1:0] __variable_wdata_961;
  assign stream_matmul_23__reduce_reset_data = __variable_wdata_961;
  reg _tmp_1525;
  reg _tmp_1526;
  reg _tmp_1527;
  reg _tmp_1528;
  assign _stream_matmul_23_source_stop = _stream_matmul_23_stream_oready && (_stream_matmul_23_source_11_idle && _stream_matmul_23_source_13_idle && _stream_matmul_23_source_15_idle && _stream_matmul_23_source_20_idle && _stream_matmul_23_source_21_idle && _stream_matmul_23_source_7_idle && _stream_matmul_23_source_9_idle && (_stream_matmul_23_fsm == 3));
  localparam _tmp_1529 = 1;
  wire [_tmp_1529-1:0] _tmp_1530;
  assign _tmp_1530 = _stream_matmul_23_source_11_idle && _stream_matmul_23_source_13_idle && _stream_matmul_23_source_15_idle && _stream_matmul_23_source_20_idle && _stream_matmul_23_source_21_idle && _stream_matmul_23_source_7_idle && _stream_matmul_23_source_9_idle && (_stream_matmul_23_fsm == 3);
  reg [_tmp_1529-1:0] _tmp_1531;
  localparam _tmp_1532 = 1;
  wire [_tmp_1532-1:0] _tmp_1533;
  assign _tmp_1533 = _stream_matmul_23_source_11_idle && _stream_matmul_23_source_13_idle && _stream_matmul_23_source_15_idle && _stream_matmul_23_source_20_idle && _stream_matmul_23_source_21_idle && _stream_matmul_23_source_7_idle && _stream_matmul_23_source_9_idle && (_stream_matmul_23_fsm == 3);
  reg [_tmp_1532-1:0] _tmp_1534;
  reg _tmp_1535;
  reg _tmp_1536;
  reg _tmp_1537;
  reg _tmp_1538;
  reg _tmp_1539;
  reg _tmp_1540;
  reg _tmp_1541;
  reg _tmp_1542;
  reg _tmp_1543;
  reg _tmp_1544;
  reg _tmp_1545;
  reg _tmp_1546;
  reg _tmp_1547;
  reg _tmp_1548;
  reg _tmp_1549;
  reg _tmp_1550;
  reg _tmp_1551;
  reg _tmp_1552;
  reg _tmp_1553;
  reg _tmp_1554;
  reg _tmp_1555;
  reg _tmp_1556;
  reg _tmp_1557;
  reg _tmp_1558;
  reg _tmp_1559;
  reg _tmp_1560;
  reg _tmp_1561;
  reg _tmp_1562;
  reg _tmp_1563;
  reg _tmp_1564;
  reg _tmp_1565;
  assign _stream_matmul_23_sink_start = _tmp_1565;
  reg _tmp_1566;
  reg _tmp_1567;
  reg _tmp_1568;
  reg _tmp_1569;
  reg _tmp_1570;
  reg _tmp_1571;
  reg _tmp_1572;
  reg _tmp_1573;
  reg _tmp_1574;
  reg _tmp_1575;
  reg _tmp_1576;
  reg _tmp_1577;
  reg _tmp_1578;
  reg _tmp_1579;
  reg _tmp_1580;
  reg _tmp_1581;
  reg _tmp_1582;
  reg _tmp_1583;
  reg _tmp_1584;
  reg _tmp_1585;
  reg _tmp_1586;
  reg _tmp_1587;
  reg _tmp_1588;
  reg _tmp_1589;
  reg _tmp_1590;
  reg _tmp_1591;
  reg _tmp_1592;
  reg _tmp_1593;
  reg _tmp_1594;
  reg _tmp_1595;
  reg _tmp_1596;
  assign _stream_matmul_23_sink_stop = _tmp_1596;
  reg _tmp_1597;
  reg _tmp_1598;
  reg _tmp_1599;
  reg _tmp_1600;
  reg _tmp_1601;
  reg _tmp_1602;
  reg _tmp_1603;
  reg _tmp_1604;
  reg _tmp_1605;
  reg _tmp_1606;
  reg _tmp_1607;
  reg _tmp_1608;
  reg _tmp_1609;
  reg _tmp_1610;
  reg _tmp_1611;
  reg _tmp_1612;
  reg _tmp_1613;
  reg _tmp_1614;
  reg _tmp_1615;
  reg _tmp_1616;
  reg _tmp_1617;
  reg _tmp_1618;
  reg _tmp_1619;
  reg _tmp_1620;
  reg _tmp_1621;
  reg _tmp_1622;
  reg _tmp_1623;
  reg _tmp_1624;
  reg _tmp_1625;
  reg _tmp_1626;
  reg _tmp_1627;
  assign _stream_matmul_23_sink_busy = _tmp_1627;
  reg _tmp_1628;
  assign _stream_matmul_23_busy = _stream_matmul_23_source_busy || _stream_matmul_23_sink_busy || _stream_matmul_23_busy_reg;
  wire matmul_23_dma_out_mask_0;
  assign matmul_23_dma_out_mask_0 = matmul_23_out_row_count + 0 >= cparam_matmul_23_out_num_row;
  wire [32-1:0] _dma_write_packed_high_local_size_1629;
  assign _dma_write_packed_high_local_size_1629 = matmul_23_next_out_write_size >> 1;
  wire [1-1:0] _dma_write_packed_low_local_size_1630;
  assign _dma_write_packed_low_local_size_1630 = matmul_23_next_out_write_size & { 1{ 1'd1 } };
  wire [32-1:0] _dma_write_packed_local_packed_size_1631;
  assign _dma_write_packed_local_packed_size_1631 = (_dma_write_packed_low_local_size_1630 > 0)? _dma_write_packed_high_local_size_1629 + 1 : _dma_write_packed_high_local_size_1629;
  wire [32-1:0] mask_addr_shifted_1632;
  assign mask_addr_shifted_1632 = matmul_23_objaddr + (matmul_23_out_base_offset + cparam_matmul_23_out_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1633;
  assign mask_addr_masked_1633 = mask_addr_shifted_1632 << 2;
  wire matmul_23_update_filter;
  assign matmul_23_update_filter = (cparam_matmul_23_data_stationary == 0) && (matmul_23_row_count >= cparam_matmul_23_max_row_count) && (matmul_23_bat_count >= cparam_matmul_23_max_bat_count) || (cparam_matmul_23_data_stationary == 1) && !cparam_matmul_23_keep_filter;
  wire matmul_23_update_act;
  assign matmul_23_update_act = (cparam_matmul_23_data_stationary == 1) && (matmul_23_och_count >= cparam_matmul_23_max_och_count) || (cparam_matmul_23_data_stationary == 0);
  wire matmul_23_mux_next_dma_flag_0;
  assign matmul_23_mux_next_dma_flag_0 = (matmul_23_row_select == 0)? (matmul_23_row_count >= cparam_matmul_23_max_row_count)? 1 : cparam_matmul_23_dma_flag_conds_0 : 1'd0;
  reg [32-1:0] matmul_33_objaddr;
  reg [32-1:0] matmul_33_arg_objaddr_0;
  reg [32-1:0] matmul_33_arg_objaddr_1;
  reg [32-1:0] matmul_33_arg_objaddr_2;
  reg [32-1:0] matmul_33_arg_objaddr_3;
  reg [32-1:0] control_matmul_33;
  localparam control_matmul_33_init = 0;
  reg _control_matmul_33_called;
  wire signed [32-1:0] matmul_33_act_base_offset;
  reg signed [32-1:0] matmul_33_act_base_offset_row;
  reg signed [32-1:0] matmul_33_act_base_offset_bat;
  assign matmul_33_act_base_offset = matmul_33_act_base_offset_row + matmul_33_act_base_offset_bat;
  reg signed [32-1:0] matmul_33_filter_base_offset;
  reg [32-1:0] matmul_33_next_stream_num_ops;
  wire signed [32-1:0] matmul_33_out_base_offset;
  reg signed [32-1:0] matmul_33_out_base_offset_val;
  reg signed [32-1:0] matmul_33_out_base_offset_col;
  reg signed [32-1:0] matmul_33_out_base_offset_row;
  reg signed [32-1:0] matmul_33_out_base_offset_bat;
  reg signed [32-1:0] matmul_33_out_base_offset_och;
  assign matmul_33_out_base_offset = matmul_33_out_base_offset_val + matmul_33_out_base_offset_col + matmul_33_out_base_offset_row + matmul_33_out_base_offset_bat + matmul_33_out_base_offset_och;
  reg matmul_33_dma_flag_0;
  reg [32-1:0] matmul_33_sync_comp_count;
  reg [32-1:0] matmul_33_sync_out_count;
  reg [32-1:0] matmul_33_write_count;
  reg [32-1:0] matmul_33_next_out_write_size;
  reg [32-1:0] matmul_33_col_count;
  reg [32-1:0] matmul_33_row_count;
  reg [32-1:0] matmul_33_bat_count;
  reg [32-1:0] matmul_33_och_count;
  reg [1-1:0] matmul_33_col_select;
  reg [1-1:0] matmul_33_row_select;
  reg [32-1:0] matmul_33_out_col_count;
  reg [32-1:0] matmul_33_out_row_count;
  reg [32-1:0] matmul_33_out_ram_select;
  reg [32-1:0] matmul_33_prev_col_count;
  reg [32-1:0] matmul_33_prev_row_count;
  reg [32-1:0] matmul_33_prev_bat_count;
  reg [32-1:0] matmul_33_prev_och_count;
  reg [1-1:0] matmul_33_prev_row_select;
  reg [32-1:0] matmul_33_stream_act_local_0;
  reg [32-1:0] matmul_33_stream_out_local_val;
  reg [32-1:0] matmul_33_stream_out_local_col;
  wire [32-1:0] matmul_33_stream_out_local;
  assign matmul_33_stream_out_local = matmul_33_stream_out_local_val + matmul_33_stream_out_local_col;
  reg [32-1:0] matmul_33_act_page_comp_offset_0;
  reg [32-1:0] matmul_33_act_page_dma_offset_0;
  reg [32-1:0] matmul_33_filter_page_comp_offset;
  reg [32-1:0] matmul_33_filter_page_dma_offset;
  reg matmul_33_out_page;
  reg [32-1:0] matmul_33_out_page_comp_offset;
  reg [32-1:0] matmul_33_out_page_dma_offset;
  reg [32-1:0] matmul_33_out_laddr_offset;
  reg matmul_33_skip_read_filter;
  reg matmul_33_skip_read_act;
  reg matmul_33_skip_comp;
  reg matmul_33_skip_write_out;
  wire [32-1:0] mask_addr_shifted_1634;
  assign mask_addr_shifted_1634 = matmul_33_arg_objaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1635;
  assign mask_addr_masked_1635 = mask_addr_shifted_1634 << 2;
  reg [32-1:0] write_burst_fsm_31;
  localparam write_burst_fsm_31_init = 0;
  reg [7-1:0] write_burst_addr_1636;
  reg [7-1:0] write_burst_stride_1637;
  reg [33-1:0] write_burst_length_1638;
  reg write_burst_done_1639;
  assign ram_w32_l128_id1_1_addr = ((write_burst_fsm_31 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_1636 : 'hx;
  assign ram_w32_l128_id1_1_wdata = ((write_burst_fsm_31 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id1_1_wenable = ((write_burst_fsm_31 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l128_id1_1_enable = ((write_burst_fsm_31 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [32-1:0] mask_addr_shifted_1640;
  assign mask_addr_shifted_1640 = matmul_33_arg_objaddr_3 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1641;
  assign mask_addr_masked_1641 = mask_addr_shifted_1640 << 2;
  reg [32-1:0] write_burst_fsm_32;
  localparam write_burst_fsm_32_init = 0;
  reg [7-1:0] write_burst_addr_1642;
  reg [7-1:0] write_burst_stride_1643;
  reg [33-1:0] write_burst_length_1644;
  reg write_burst_done_1645;
  assign ram_w32_l128_id2_1_addr = ((write_burst_fsm_32 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_1642 : 'hx;
  assign ram_w32_l128_id2_1_wdata = ((write_burst_fsm_32 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id2_1_wenable = ((write_burst_fsm_32 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l128_id2_1_enable = ((write_burst_fsm_32 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [32-1:0] mask_addr_shifted_1646;
  assign mask_addr_shifted_1646 = matmul_33_arg_objaddr_1 + matmul_33_filter_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1647;
  assign mask_addr_masked_1647 = mask_addr_shifted_1646 << 2;
  wire write_burst_block_ram_wvalid_1648;
  wire write_burst_block_ram_wquit_1649;
  reg [32-1:0] write_burst_fsm_33;
  localparam write_burst_fsm_33_init = 0;
  reg [9-1:0] write_burst_addr_1650;
  reg [9-1:0] write_burst_stride_1651;
  reg [33-1:0] write_burst_length_1652;
  reg write_burst_done_1653;
  assign ram_w32_l512_id1_1_addr = ((write_burst_fsm_33 == 1) && write_burst_block_ram_wvalid_1648)? write_burst_addr_1650 : 'hx;
  assign ram_w32_l512_id1_1_wdata = ((write_burst_fsm_33 == 1) && write_burst_block_ram_wvalid_1648)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l512_id1_1_wenable = ((write_burst_fsm_33 == 1) && write_burst_block_ram_wvalid_1648)? 1'd1 : 0;
  assign ram_w32_l512_id1_1_enable = ((write_burst_fsm_33 == 1) && write_burst_block_ram_wvalid_1648)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_1654;
  wire write_burst_block_ram_wquit_1655;
  reg [32-1:0] write_burst_fsm_34;
  localparam write_burst_fsm_34_init = 0;
  reg [10-1:0] write_burst_addr_1656;
  reg [10-1:0] write_burst_stride_1657;
  reg [33-1:0] write_burst_length_1658;
  reg write_burst_done_1659;
  assign ram_w32_l1024_id0_1_addr = ((write_burst_fsm_34 == 1) && write_burst_block_ram_wvalid_1654)? write_burst_addr_1656 : 
                                    ((read_burst_fsm_26 == 1) && (!read_burst_rvalid_1301 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_addr_1298 : 'hx;
  assign ram_w32_l1024_id0_1_wdata = ((write_burst_fsm_34 == 1) && write_burst_block_ram_wvalid_1654)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l1024_id0_1_wenable = ((write_burst_fsm_34 == 1) && write_burst_block_ram_wvalid_1654)? 1'd1 : 0;
  assign ram_w32_l1024_id0_1_enable = ((write_burst_fsm_34 == 1) && write_burst_block_ram_wvalid_1654)? 1'd1 : 
                                      ((read_burst_fsm_26 == 1) && (!read_burst_rvalid_1301 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_35;
  localparam write_burst_block_fsm_35_init = 0;
  reg [33-1:0] write_burst_block_length_1660;
  reg [32-1:0] write_burst_block_blocksize_1661;
  reg write_burst_block_done_1662;
  reg [32-1:0] write_burst_block_count_1663;
  assign write_burst_block_ram_wvalid_1648 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_35 == 1);
  assign write_burst_block_ram_wquit_1649 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_1660 <= 1);
  assign write_burst_block_ram_wvalid_1654 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_35 == 2);
  assign write_burst_block_ram_wquit_1655 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_1660 <= 1);
  wire [32-1:0] matmul_33_mux_act_gaddr_0;
  assign matmul_33_mux_act_gaddr_0 = (matmul_33_row_select == 0)? matmul_33_arg_objaddr_0 + (matmul_33_act_base_offset + cparam_matmul_33_act_offset_values_0) : 1'd0;
  wire matmul_33_dma_pad_mask_0;
  assign matmul_33_dma_pad_mask_0 = (matmul_33_row_count + 0 < cparam_matmul_33_pad_row_top) || (matmul_33_row_count + 0 >= cparam_matmul_33_act_num_row + cparam_matmul_33_pad_row_top);
  wire matmul_33_mux_dma_pad_mask_0;
  assign matmul_33_mux_dma_pad_mask_0 = (matmul_33_row_select == 0)? matmul_33_dma_pad_mask_0 : 1'd0;
  wire matmul_33_mux_dma_flag_0;
  assign matmul_33_mux_dma_flag_0 = (matmul_33_prev_row_select == 0)? matmul_33_dma_flag_0 : 1'd0;
  wire [32-1:0] mask_addr_shifted_1664;
  assign mask_addr_shifted_1664 = matmul_33_mux_act_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1665;
  assign mask_addr_masked_1665 = mask_addr_shifted_1664 << 2;
  assign _maxi_read_req_fifo_deq = ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 15)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 14)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 13)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 12)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 11)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 10)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1)) && !_maxi_read_req_fifo_empty)? 1 : 0;
  reg [32-1:0] write_burst_fsm_36;
  localparam write_burst_fsm_36_init = 0;
  reg [9-1:0] write_burst_addr_1666;
  reg [9-1:0] write_burst_stride_1667;
  reg [33-1:0] write_burst_length_1668;
  reg write_burst_done_1669;
  assign ram_w32_l512_id0_1_addr = ((write_burst_fsm_36 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_1666 : 'hx;
  assign ram_w32_l512_id0_1_wdata = ((write_burst_fsm_36 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l512_id0_1_wenable = ((write_burst_fsm_36 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l512_id0_1_enable = ((write_burst_fsm_36 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign _maxi_rready_sb_0 = (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2);
  reg [32-1:0] matmul_33_comp_fsm;
  localparam matmul_33_comp_fsm_init = 0;
  reg [32-1:0] matmul_33_filter_page_comp_offset_buf;
  reg [32-1:0] matmul_33_act_page_comp_offset_buf_0;
  reg [32-1:0] matmul_33_out_page_comp_offset_buf;
  reg [32-1:0] matmul_33_row_count_buf;
  reg [1-1:0] matmul_33_row_select_buf;
  reg [32-1:0] matmul_33_och_count_buf;
  wire matmul_33_stream_pad_mask_0_0;
  assign matmul_33_stream_pad_mask_0_0 = (matmul_33_col_count + 0 < cparam_matmul_33_pad_col_left) || (matmul_33_col_count + 0 >= cparam_matmul_33_act_num_col + cparam_matmul_33_pad_col_left) || (matmul_33_row_count_buf + 0 < cparam_matmul_33_pad_row_top) || (matmul_33_row_count_buf + 0 >= cparam_matmul_33_act_num_row + cparam_matmul_33_pad_row_top);
  reg [1-1:0] matmul_33_stream_pad_masks;
  wire [9-1:0] stream_matmul_33_parameter_0_data;
  wire [1-1:0] stream_matmul_33_parameter_1_data;
  wire [1-1:0] stream_matmul_33_parameter_2_data;
  wire [1-1:0] stream_matmul_33_parameter_3_data;
  wire [2-1:0] stream_matmul_33_parameter_4_data;
  wire [1-1:0] stream_matmul_33__reduce_reset_data;
  wire [1-1:0] stream_matmul_33_parameter_6_data;
  wire [32-1:0] stream_matmul_33_source_7_data;
  wire [1-1:0] stream_matmul_33_parameter_8_data;
  wire [32-1:0] stream_matmul_33_source_9_data;
  wire [1-1:0] stream_matmul_33_parameter_10_data;
  wire [32-1:0] stream_matmul_33_source_11_data;
  wire [1-1:0] stream_matmul_33_parameter_12_data;
  wire [32-1:0] stream_matmul_33_source_13_data;
  wire [1-1:0] stream_matmul_33_parameter_14_data;
  wire [32-1:0] stream_matmul_33_source_15_data;
  wire [1-1:0] stream_matmul_33_parameter_16_data;
  wire [1-1:0] stream_matmul_33_parameter_17_data;
  wire [5-1:0] stream_matmul_33_parameter_18_data;
  wire [1-1:0] stream_matmul_33_parameter_19_data;
  wire [32-1:0] stream_matmul_33_source_20_data;
  wire [32-1:0] stream_matmul_33_source_21_data;
  wire [32-1:0] stream_matmul_33_source_22_data;
  reg __stream_matmul_33_stream_ivalid_1;
  reg __stream_matmul_33_stream_ivalid_2;
  reg __stream_matmul_33_stream_ivalid_3;
  reg __stream_matmul_33_stream_ivalid_4;
  reg __stream_matmul_33_stream_ivalid_5;
  reg __stream_matmul_33_stream_ivalid_6;
  reg __stream_matmul_33_stream_ivalid_7;
  reg __stream_matmul_33_stream_ivalid_8;
  reg __stream_matmul_33_stream_ivalid_9;
  reg __stream_matmul_33_stream_ivalid_10;
  reg __stream_matmul_33_stream_ivalid_11;
  reg __stream_matmul_33_stream_ivalid_12;
  reg __stream_matmul_33_stream_ivalid_13;
  reg __stream_matmul_33_stream_ivalid_14;
  reg __stream_matmul_33_stream_ivalid_15;
  reg __stream_matmul_33_stream_ivalid_16;
  reg __stream_matmul_33_stream_ivalid_17;
  reg __stream_matmul_33_stream_ivalid_18;
  reg __stream_matmul_33_stream_ivalid_19;
  reg __stream_matmul_33_stream_ivalid_20;
  reg __stream_matmul_33_stream_ivalid_21;
  reg __stream_matmul_33_stream_ivalid_22;
  reg __stream_matmul_33_stream_ivalid_23;
  reg __stream_matmul_33_stream_ivalid_24;
  reg __stream_matmul_33_stream_ivalid_25;
  reg __stream_matmul_33_stream_ivalid_26;
  reg __stream_matmul_33_stream_ivalid_27;
  reg __stream_matmul_33_stream_ivalid_28;
  reg __stream_matmul_33_stream_ivalid_29;
  reg __stream_matmul_33_stream_ivalid_30;
  reg [32-1:0] _counter_data_1058;
  reg [32-1:0] _counter_count_1058;
  wire _counter_reset_cond_1058;
  assign _counter_reset_cond_1058 = stream_matmul_33__reduce_reset_data;
  wire [32-1:0] _counter_current_count_1058;
  assign _counter_current_count_1058 = (_counter_reset_cond_1058)? 1'sd0 : _counter_count_1058;
  wire [1-1:0] _pointer_data_1061;
  assign _pointer_data_1061 = stream_matmul_33_parameter_4_data[1'sd0];
  reg [9-1:0] _minus_data_1063;
  wire [1-1:0] _pointer_data_1067;
  assign _pointer_data_1067 = stream_matmul_33_parameter_4_data[2'sd1];
  reg [9-1:0] _minus_data_1069;
  wire [16-1:0] _slice_data_1077;
  assign _slice_data_1077 = stream_matmul_33_source_7_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1078;
  assign _reinterpretcast_src_1078 = _slice_data_1077;
  wire signed [16-1:0] _reinterpretcast_data_1078;
  assign _reinterpretcast_data_1078 = _reinterpretcast_src_1078;
  wire [16-1:0] _slice_data_1081;
  assign _slice_data_1081 = stream_matmul_33_source_7_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1082;
  assign _reinterpretcast_src_1082 = _slice_data_1081;
  wire signed [16-1:0] _reinterpretcast_data_1082;
  assign _reinterpretcast_data_1082 = _reinterpretcast_src_1082;
  wire signed [16-1:0] _cond_data_1083;
  assign _cond_data_1083 = (stream_matmul_33_parameter_6_data)? _reinterpretcast_data_1078 : _reinterpretcast_data_1078;
  wire signed [16-1:0] _cond_data_1084;
  assign _cond_data_1084 = (stream_matmul_33_parameter_6_data)? _reinterpretcast_data_1078 : _reinterpretcast_data_1082;
  wire [16-1:0] _slice_data_1089;
  assign _slice_data_1089 = stream_matmul_33_source_9_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1090;
  assign _reinterpretcast_src_1090 = _slice_data_1089;
  wire signed [16-1:0] _reinterpretcast_data_1090;
  assign _reinterpretcast_data_1090 = _reinterpretcast_src_1090;
  wire [16-1:0] _slice_data_1093;
  assign _slice_data_1093 = stream_matmul_33_source_9_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1094;
  assign _reinterpretcast_src_1094 = _slice_data_1093;
  wire signed [16-1:0] _reinterpretcast_data_1094;
  assign _reinterpretcast_data_1094 = _reinterpretcast_src_1094;
  wire signed [16-1:0] _cond_data_1095;
  assign _cond_data_1095 = (stream_matmul_33_parameter_8_data)? _reinterpretcast_data_1090 : _reinterpretcast_data_1090;
  wire signed [16-1:0] _cond_data_1096;
  assign _cond_data_1096 = (stream_matmul_33_parameter_8_data)? _reinterpretcast_data_1090 : _reinterpretcast_data_1094;
  wire [16-1:0] _slice_data_1101;
  assign _slice_data_1101 = stream_matmul_33_source_11_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1102;
  assign _reinterpretcast_src_1102 = _slice_data_1101;
  wire [16-1:0] _reinterpretcast_data_1102;
  assign _reinterpretcast_data_1102 = _reinterpretcast_src_1102;
  wire [16-1:0] _slice_data_1105;
  assign _slice_data_1105 = stream_matmul_33_source_11_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1106;
  assign _reinterpretcast_src_1106 = _slice_data_1105;
  wire [16-1:0] _reinterpretcast_data_1106;
  assign _reinterpretcast_data_1106 = _reinterpretcast_src_1106;
  wire [16-1:0] _cond_data_1107;
  assign _cond_data_1107 = (stream_matmul_33_parameter_10_data)? _reinterpretcast_data_1102 : _reinterpretcast_data_1102;
  wire [16-1:0] _cond_data_1108;
  assign _cond_data_1108 = (stream_matmul_33_parameter_10_data)? _reinterpretcast_data_1102 : _reinterpretcast_data_1106;
  wire [16-1:0] _slice_data_1113;
  assign _slice_data_1113 = stream_matmul_33_source_13_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1114;
  assign _reinterpretcast_src_1114 = _slice_data_1113;
  wire [16-1:0] _reinterpretcast_data_1114;
  assign _reinterpretcast_data_1114 = _reinterpretcast_src_1114;
  wire [16-1:0] _slice_data_1117;
  assign _slice_data_1117 = stream_matmul_33_source_13_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1118;
  assign _reinterpretcast_src_1118 = _slice_data_1117;
  wire [16-1:0] _reinterpretcast_data_1118;
  assign _reinterpretcast_data_1118 = _reinterpretcast_src_1118;
  wire [16-1:0] _cond_data_1119;
  assign _cond_data_1119 = (stream_matmul_33_parameter_12_data)? _reinterpretcast_data_1114 : _reinterpretcast_data_1114;
  wire [16-1:0] _cond_data_1120;
  assign _cond_data_1120 = (stream_matmul_33_parameter_12_data)? _reinterpretcast_data_1114 : _reinterpretcast_data_1118;
  wire [16-1:0] _slice_data_1125;
  assign _slice_data_1125 = stream_matmul_33_source_15_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1126;
  assign _reinterpretcast_src_1126 = _slice_data_1125;
  wire [16-1:0] _reinterpretcast_data_1126;
  assign _reinterpretcast_data_1126 = _reinterpretcast_src_1126;
  wire [16-1:0] _slice_data_1129;
  assign _slice_data_1129 = stream_matmul_33_source_15_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1130;
  assign _reinterpretcast_src_1130 = _slice_data_1129;
  wire [16-1:0] _reinterpretcast_data_1130;
  assign _reinterpretcast_data_1130 = _reinterpretcast_src_1130;
  wire [16-1:0] _cond_data_1131;
  assign _cond_data_1131 = (stream_matmul_33_parameter_14_data)? _reinterpretcast_data_1126 : _reinterpretcast_data_1126;
  wire [16-1:0] _cond_data_1132;
  assign _cond_data_1132 = (stream_matmul_33_parameter_14_data)? _reinterpretcast_data_1126 : _reinterpretcast_data_1130;
  reg [1-1:0] _eq_data_1138;
  reg [1-1:0] _eq_data_1142;
  wire [16-1:0] _slice_data_1162;
  assign _slice_data_1162 = stream_matmul_33_source_21_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1163;
  assign _reinterpretcast_src_1163 = _slice_data_1162;
  wire signed [16-1:0] _reinterpretcast_data_1163;
  assign _reinterpretcast_data_1163 = _reinterpretcast_src_1163;
  wire [16-1:0] _slice_data_1166;
  assign _slice_data_1166 = stream_matmul_33_source_21_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1167;
  assign _reinterpretcast_src_1167 = _slice_data_1166;
  wire signed [16-1:0] _reinterpretcast_data_1167;
  assign _reinterpretcast_data_1167 = _reinterpretcast_src_1167;
  wire [16-1:0] _slice_data_1174;
  assign _slice_data_1174 = stream_matmul_33_source_22_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1175;
  assign _reinterpretcast_src_1175 = _slice_data_1174;
  wire signed [16-1:0] _reinterpretcast_data_1175;
  assign _reinterpretcast_data_1175 = _reinterpretcast_src_1175;
  wire [16-1:0] _slice_data_1178;
  assign _slice_data_1178 = stream_matmul_33_source_22_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1179;
  assign _reinterpretcast_src_1179 = _slice_data_1178;
  wire signed [16-1:0] _reinterpretcast_data_1179;
  assign _reinterpretcast_data_1179 = _reinterpretcast_src_1179;
  wire [1-1:0] _pointer_data_1184;
  assign _pointer_data_1184 = stream_matmul_33_parameter_3_data[1'sd0];
  reg [16-1:0] _plus_data_1189;
  reg [16-1:0] _plus_data_1194;
  reg [16-1:0] _plus_data_1199;
  reg [16-1:0] _plus_data_1204;
  reg [16-1:0] _plus_data_1210;
  reg [16-1:0] _plus_data_1215;
  reg [16-1:0] _plus_data_1231;
  reg [16-1:0] _plus_data_1250;
  reg [1-1:0] __delay_data_1501_pointer_1061;
  reg [32-1:0] __delay_data_1503__variable_1137;
  reg [1-1:0] __delay_data_1506_pointer_1184;
  reg signed [16-1:0] __delay_data_1509_reinterpretcast_1163;
  reg [1-1:0] __delay_data_1514_pointer_1067;
  reg signed [16-1:0] __delay_data_1518_reinterpretcast_1167;
  reg [1-1:0] __delay_data_1523__variable_1057;
  reg [9-1:0] __delay_data_1550__variable_1052;
  reg signed [16-1:0] __delay_data_1564_reinterpretcast_1175;
  reg signed [16-1:0] __delay_data_1569_reinterpretcast_1179;
  reg signed [16-1:0] __delay_data_1587_cond_1084;
  reg signed [16-1:0] __delay_data_1607_cond_1096;
  reg signed [16-1:0] __delay_data_1648_cond_1083;
  reg signed [16-1:0] __delay_data_1668_cond_1095;
  reg [1-1:0] _eq_data_1065;
  reg [1-1:0] _eq_data_1071;
  wire signed [32-1:0] _cond_data_1140;
  assign _cond_data_1140 = (_eq_data_1138)? __delay_data_1503__variable_1137 : 1'sd0;
  wire signed [32-1:0] _cond_data_1144;
  assign _cond_data_1144 = (_eq_data_1142)? _cond_data_1140 : 1'sd0;
  wire [16-1:0] _slice_data_1148;
  assign _slice_data_1148 = _cond_data_1144[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1149;
  assign _reinterpretcast_src_1149 = _slice_data_1148;
  wire signed [16-1:0] _reinterpretcast_data_1149;
  assign _reinterpretcast_data_1149 = _reinterpretcast_src_1149;
  wire [16-1:0] _slice_data_1152;
  assign _slice_data_1152 = _cond_data_1144[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1153;
  assign _reinterpretcast_src_1153 = _slice_data_1152;
  wire signed [16-1:0] _reinterpretcast_data_1153;
  assign _reinterpretcast_data_1153 = _reinterpretcast_src_1153;
  reg [1-1:0] __delay_data_1502__delay_1501_pointer_1061;
  reg signed [16-1:0] __delay_data_1504_reinterpretcast_1149;
  reg [1-1:0] __delay_data_1507__delay_1506_pointer_1184;
  reg signed [16-1:0] __delay_data_1510__delay_1509_reinterpretcast_1163;
  reg [16-1:0] __delay_data_1512_plus_1189;
  reg [1-1:0] __delay_data_1515__delay_1514_pointer_1067;
  reg signed [16-1:0] __delay_data_1516_reinterpretcast_1153;
  reg signed [16-1:0] __delay_data_1519__delay_1518_reinterpretcast_1167;
  reg [16-1:0] __delay_data_1521_plus_1194;
  reg [1-1:0] __delay_data_1524__delay_1523__variable_1057;
  reg [16-1:0] __delay_data_1537_plus_1199;
  reg [9-1:0] __delay_data_1551__delay_1550__variable_1052;
  reg signed [16-1:0] __delay_data_1565__delay_1564_reinterpretcast_1175;
  reg [16-1:0] __delay_data_1567_plus_1210;
  reg signed [16-1:0] __delay_data_1570__delay_1569_reinterpretcast_1179;
  reg [16-1:0] __delay_data_1572_plus_1215;
  reg [16-1:0] __delay_data_1574_plus_1231;
  reg signed [16-1:0] __delay_data_1588__delay_1587_cond_1084;
  reg signed [16-1:0] __delay_data_1608__delay_1607_cond_1096;
  reg [16-1:0] __delay_data_1628_plus_1250;
  reg signed [16-1:0] __delay_data_1649__delay_1648_cond_1083;
  reg signed [16-1:0] __delay_data_1669__delay_1668_cond_1095;
  reg [16-1:0] __delay_data_1689_plus_1204;
  reg [1-1:0] _land_data_1066;
  reg [1-1:0] _land_data_1072;
  reg signed [16-1:0] __delay_data_1505__delay_1504_reinterpretcast_1149;
  reg [1-1:0] __delay_data_1508__delay_1507__delay_1506_pointer_1184;
  reg signed [16-1:0] __delay_data_1511__delay_1510__delay_1509_reinterpretcast_1163;
  reg [16-1:0] __delay_data_1513__delay_1512_plus_1189;
  reg signed [16-1:0] __delay_data_1517__delay_1516_reinterpretcast_1153;
  reg signed [16-1:0] __delay_data_1520__delay_1519__delay_1518_reinterpretcast_1167;
  reg [16-1:0] __delay_data_1522__delay_1521_plus_1194;
  reg [1-1:0] __delay_data_1525__delay_1524__delay_1523__variable_1057;
  reg [16-1:0] __delay_data_1538__delay_1537_plus_1199;
  reg [9-1:0] __delay_data_1552__delay_1551__delay_1550__variable_1052;
  reg signed [16-1:0] __delay_data_1566__delay_1565__delay_1564_reinterpretcast_1175;
  reg [16-1:0] __delay_data_1568__delay_1567_plus_1210;
  reg signed [16-1:0] __delay_data_1571__delay_1570__delay_1569_reinterpretcast_1179;
  reg [16-1:0] __delay_data_1573__delay_1572_plus_1215;
  reg [16-1:0] __delay_data_1575__delay_1574_plus_1231;
  reg signed [16-1:0] __delay_data_1589__delay_1588__delay_1587_cond_1084;
  reg signed [16-1:0] __delay_data_1609__delay_1608__delay_1607_cond_1096;
  reg [16-1:0] __delay_data_1629__delay_1628_plus_1250;
  reg signed [16-1:0] __delay_data_1650__delay_1649__delay_1648_cond_1083;
  reg signed [16-1:0] __delay_data_1670__delay_1669__delay_1668_cond_1095;
  reg [16-1:0] __delay_data_1690__delay_1689_plus_1204;
  wire signed [16-1:0] _cond_data_1155;
  assign _cond_data_1155 = (_land_data_1066)? 1'sd0 : __delay_data_1505__delay_1504_reinterpretcast_1149;
  wire signed [16-1:0] _cond_data_1157;
  assign _cond_data_1157 = (_land_data_1072)? 1'sd0 : __delay_data_1517__delay_1516_reinterpretcast_1153;
  wire signed [16-1:0] _cond_data_1169;
  assign _cond_data_1169 = (_land_data_1066)? 1'sd0 : __delay_data_1511__delay_1510__delay_1509_reinterpretcast_1163;
  wire signed [16-1:0] _cond_data_1171;
  assign _cond_data_1171 = (_land_data_1072)? 1'sd0 : __delay_data_1520__delay_1519__delay_1518_reinterpretcast_1167;
  wire signed [16-1:0] _cond_data_1181;
  assign _cond_data_1181 = (_land_data_1066)? 1'sd0 : __delay_data_1566__delay_1565__delay_1564_reinterpretcast_1175;
  wire signed [16-1:0] _cond_data_1183;
  assign _cond_data_1183 = (_land_data_1072)? 1'sd0 : __delay_data_1571__delay_1570__delay_1569_reinterpretcast_1179;
  wire signed [16-1:0] _cond_data_1187;
  assign _cond_data_1187 = (__delay_data_1508__delay_1507__delay_1506_pointer_1184)? 1'sd0 : _cond_data_1155;
  assign _mul_8_is_root = ((_stream_matmul_33_busy)? 0 : 1) && (((_stream_matmul_23_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1));
  assign _mul_8_stream_oready = ((_stream_matmul_33_busy)? _stream_matmul_33_stream_oready : 1) && (((_stream_matmul_23_busy)? _stream_matmul_23_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_8_stream_internal_oready));
  wire signed [16-1:0] _cond_data_1192;
  assign _cond_data_1192 = (__delay_data_1508__delay_1507__delay_1506_pointer_1184)? 1'sd0 : _cond_data_1157;
  assign _mul_9_is_root = ((_stream_matmul_33_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _mul_9_stream_oready = ((_stream_matmul_33_busy)? _stream_matmul_33_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_9_stream_internal_oready);
  wire signed [16-1:0] _cond_data_1208;
  assign _cond_data_1208 = (__delay_data_1508__delay_1507__delay_1506_pointer_1184)? 1'sd0 : _cond_data_1155;
  assign _mul_10_is_root = ((_stream_matmul_33_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _mul_10_stream_oready = ((_stream_matmul_33_busy)? _stream_matmul_33_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_10_stream_internal_oready);
  wire signed [16-1:0] _cond_data_1213;
  assign _cond_data_1213 = (__delay_data_1508__delay_1507__delay_1506_pointer_1184)? 1'sd0 : _cond_data_1157;
  assign _mul_11_is_root = ((_stream_matmul_33_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _mul_11_stream_oready = ((_stream_matmul_33_busy)? _stream_matmul_33_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_11_stream_internal_oready);
  reg [1-1:0] __delay_data_1526__delay_1525__delay_1524____variable_1057;
  reg [16-1:0] __delay_data_1539__delay_1538__delay_1537_plus_1199;
  reg [9-1:0] __delay_data_1553__delay_1552__delay_1551____variable_1052;
  reg [16-1:0] __delay_data_1576__delay_1575__delay_1574_plus_1231;
  reg signed [16-1:0] __delay_data_1590__delay_1589__delay_1588___cond_1084;
  reg signed [16-1:0] __delay_data_1610__delay_1609__delay_1608___cond_1096;
  reg [16-1:0] __delay_data_1630__delay_1629__delay_1628_plus_1250;
  reg signed [16-1:0] __delay_data_1651__delay_1650__delay_1649___cond_1083;
  reg signed [16-1:0] __delay_data_1671__delay_1670__delay_1669___cond_1095;
  reg [16-1:0] __delay_data_1691__delay_1690__delay_1689_plus_1204;
  reg [1-1:0] __delay_data_1527__delay_1526__delay_1525____variable_1057;
  reg [16-1:0] __delay_data_1540__delay_1539__delay_1538___plus_1199;
  reg [9-1:0] __delay_data_1554__delay_1553__delay_1552____variable_1052;
  reg [16-1:0] __delay_data_1577__delay_1576__delay_1575___plus_1231;
  reg signed [16-1:0] __delay_data_1591__delay_1590__delay_1589___cond_1084;
  reg signed [16-1:0] __delay_data_1611__delay_1610__delay_1609___cond_1096;
  reg [16-1:0] __delay_data_1631__delay_1630__delay_1629___plus_1250;
  reg signed [16-1:0] __delay_data_1652__delay_1651__delay_1650___cond_1083;
  reg signed [16-1:0] __delay_data_1672__delay_1671__delay_1670___cond_1095;
  reg [16-1:0] __delay_data_1692__delay_1691__delay_1690___plus_1204;
  reg [1-1:0] __delay_data_1528__delay_1527__delay_1526____variable_1057;
  reg [16-1:0] __delay_data_1541__delay_1540__delay_1539___plus_1199;
  reg [9-1:0] __delay_data_1555__delay_1554__delay_1553____variable_1052;
  reg [16-1:0] __delay_data_1578__delay_1577__delay_1576___plus_1231;
  reg signed [16-1:0] __delay_data_1592__delay_1591__delay_1590___cond_1084;
  reg signed [16-1:0] __delay_data_1612__delay_1611__delay_1610___cond_1096;
  reg [16-1:0] __delay_data_1632__delay_1631__delay_1630___plus_1250;
  reg signed [16-1:0] __delay_data_1653__delay_1652__delay_1651___cond_1083;
  reg signed [16-1:0] __delay_data_1673__delay_1672__delay_1671___cond_1095;
  reg [16-1:0] __delay_data_1693__delay_1692__delay_1691___plus_1204;
  reg [1-1:0] __delay_data_1529__delay_1528__delay_1527____variable_1057;
  reg [16-1:0] __delay_data_1542__delay_1541__delay_1540___plus_1199;
  reg [9-1:0] __delay_data_1556__delay_1555__delay_1554____variable_1052;
  reg [16-1:0] __delay_data_1579__delay_1578__delay_1577___plus_1231;
  reg signed [16-1:0] __delay_data_1593__delay_1592__delay_1591___cond_1084;
  reg signed [16-1:0] __delay_data_1613__delay_1612__delay_1611___cond_1096;
  reg [16-1:0] __delay_data_1633__delay_1632__delay_1631___plus_1250;
  reg signed [16-1:0] __delay_data_1654__delay_1653__delay_1652___cond_1083;
  reg signed [16-1:0] __delay_data_1674__delay_1673__delay_1672___cond_1095;
  reg [16-1:0] __delay_data_1694__delay_1693__delay_1692___plus_1204;
  reg [1-1:0] __delay_data_1530__delay_1529__delay_1528____variable_1057;
  reg [16-1:0] __delay_data_1543__delay_1542__delay_1541___plus_1199;
  reg [9-1:0] __delay_data_1557__delay_1556__delay_1555____variable_1052;
  reg [16-1:0] __delay_data_1580__delay_1579__delay_1578___plus_1231;
  reg signed [16-1:0] __delay_data_1594__delay_1593__delay_1592___cond_1084;
  reg signed [16-1:0] __delay_data_1614__delay_1613__delay_1612___cond_1096;
  reg [16-1:0] __delay_data_1634__delay_1633__delay_1632___plus_1250;
  reg signed [16-1:0] __delay_data_1655__delay_1654__delay_1653___cond_1083;
  reg signed [16-1:0] __delay_data_1675__delay_1674__delay_1673___cond_1095;
  reg [16-1:0] __delay_data_1695__delay_1694__delay_1693___plus_1204;
  reg [1-1:0] __delay_data_1531__delay_1530__delay_1529____variable_1057;
  reg [16-1:0] __delay_data_1544__delay_1543__delay_1542___plus_1199;
  reg [9-1:0] __delay_data_1558__delay_1557__delay_1556____variable_1052;
  reg [16-1:0] __delay_data_1581__delay_1580__delay_1579___plus_1231;
  reg signed [16-1:0] __delay_data_1595__delay_1594__delay_1593___cond_1084;
  reg signed [16-1:0] __delay_data_1615__delay_1614__delay_1613___cond_1096;
  reg [16-1:0] __delay_data_1635__delay_1634__delay_1633___plus_1250;
  reg signed [16-1:0] __delay_data_1656__delay_1655__delay_1654___cond_1083;
  reg signed [16-1:0] __delay_data_1676__delay_1675__delay_1674___cond_1095;
  reg [16-1:0] __delay_data_1696__delay_1695__delay_1694___plus_1204;
  reg [1-1:0] __delay_data_1532__delay_1531__delay_1530____variable_1057;
  reg [16-1:0] __delay_data_1545__delay_1544__delay_1543___plus_1199;
  reg [9-1:0] __delay_data_1559__delay_1558__delay_1557____variable_1052;
  reg [16-1:0] __delay_data_1582__delay_1581__delay_1580___plus_1231;
  reg signed [16-1:0] __delay_data_1596__delay_1595__delay_1594___cond_1084;
  reg signed [16-1:0] __delay_data_1616__delay_1615__delay_1614___cond_1096;
  reg [16-1:0] __delay_data_1636__delay_1635__delay_1634___plus_1250;
  reg signed [16-1:0] __delay_data_1657__delay_1656__delay_1655___cond_1083;
  reg signed [16-1:0] __delay_data_1677__delay_1676__delay_1675___cond_1095;
  reg [16-1:0] __delay_data_1697__delay_1696__delay_1695___plus_1204;
  reg [1-1:0] __delay_data_1533__delay_1532__delay_1531____variable_1057;
  reg [16-1:0] __delay_data_1546__delay_1545__delay_1544___plus_1199;
  reg [9-1:0] __delay_data_1560__delay_1559__delay_1558____variable_1052;
  reg [16-1:0] __delay_data_1583__delay_1582__delay_1581___plus_1231;
  reg signed [16-1:0] __delay_data_1597__delay_1596__delay_1595___cond_1084;
  reg signed [16-1:0] __delay_data_1617__delay_1616__delay_1615___cond_1096;
  reg [16-1:0] __delay_data_1637__delay_1636__delay_1635___plus_1250;
  reg signed [16-1:0] __delay_data_1658__delay_1657__delay_1656___cond_1083;
  reg signed [16-1:0] __delay_data_1678__delay_1677__delay_1676___cond_1095;
  reg [16-1:0] __delay_data_1698__delay_1697__delay_1696___plus_1204;
  reg [1-1:0] __delay_data_1534__delay_1533__delay_1532____variable_1057;
  reg [16-1:0] __delay_data_1547__delay_1546__delay_1545___plus_1199;
  reg [9-1:0] __delay_data_1561__delay_1560__delay_1559____variable_1052;
  reg [16-1:0] __delay_data_1584__delay_1583__delay_1582___plus_1231;
  reg signed [16-1:0] __delay_data_1598__delay_1597__delay_1596___cond_1084;
  reg signed [16-1:0] __delay_data_1618__delay_1617__delay_1616___cond_1096;
  reg [16-1:0] __delay_data_1638__delay_1637__delay_1636___plus_1250;
  reg signed [16-1:0] __delay_data_1659__delay_1658__delay_1657___cond_1083;
  reg signed [16-1:0] __delay_data_1679__delay_1678__delay_1677___cond_1095;
  reg [16-1:0] __delay_data_1699__delay_1698__delay_1697___plus_1204;
  wire signed [32-1:0] __substreamoutput_data_1190;
  assign __substreamoutput_data_1190 = mul_8_z_data;
  wire signed [32-1:0] __substreamoutput_data_1195;
  assign __substreamoutput_data_1195 = mul_9_z_data;
  reg signed [64-1:0] __variable_wdata_46;
  assign add_tree_3_var0_data = __variable_wdata_46;
  reg signed [64-1:0] __variable_wdata_47;
  assign add_tree_3_var1_data = __variable_wdata_47;
  assign _add_tree_3_is_root = ((_stream_matmul_33_busy)? 0 : 1) && 1;
  assign _add_tree_3_stream_oready = ((_stream_matmul_33_busy)? _stream_matmul_33_stream_oready : 1) && _add_tree_3_stream_internal_oready;
  wire signed [32-1:0] __substreamoutput_data_1211;
  assign __substreamoutput_data_1211 = mul_10_z_data;
  wire signed [32-1:0] __substreamoutput_data_1216;
  assign __substreamoutput_data_1216 = mul_11_z_data;
  reg signed [64-1:0] __variable_wdata_50;
  assign add_tree_4_var0_data = __variable_wdata_50;
  reg signed [64-1:0] __variable_wdata_51;
  assign add_tree_4_var1_data = __variable_wdata_51;
  assign _add_tree_4_is_root = ((_stream_matmul_33_busy)? 0 : 1) && 1;
  assign _add_tree_4_stream_oready = ((_stream_matmul_33_busy)? _stream_matmul_33_stream_oready : 1) && _add_tree_4_stream_internal_oready;
  reg [1-1:0] __delay_data_1535__delay_1534__delay_1533____variable_1057;
  reg [16-1:0] __delay_data_1548__delay_1547__delay_1546___plus_1199;
  reg [9-1:0] __delay_data_1562__delay_1561__delay_1560____variable_1052;
  reg [16-1:0] __delay_data_1585__delay_1584__delay_1583___plus_1231;
  reg signed [16-1:0] __delay_data_1599__delay_1598__delay_1597___cond_1084;
  reg signed [16-1:0] __delay_data_1619__delay_1618__delay_1617___cond_1096;
  reg [16-1:0] __delay_data_1639__delay_1638__delay_1637___plus_1250;
  reg signed [16-1:0] __delay_data_1660__delay_1659__delay_1658___cond_1083;
  reg signed [16-1:0] __delay_data_1680__delay_1679__delay_1678___cond_1095;
  reg [16-1:0] __delay_data_1700__delay_1699__delay_1698___plus_1204;
  reg [1-1:0] __delay_data_1536__delay_1535__delay_1534____variable_1057;
  reg [16-1:0] __delay_data_1549__delay_1548__delay_1547___plus_1199;
  reg [9-1:0] __delay_data_1563__delay_1562__delay_1561____variable_1052;
  reg [16-1:0] __delay_data_1586__delay_1585__delay_1584___plus_1231;
  reg signed [16-1:0] __delay_data_1600__delay_1599__delay_1598___cond_1084;
  reg signed [16-1:0] __delay_data_1620__delay_1619__delay_1618___cond_1096;
  reg [16-1:0] __delay_data_1640__delay_1639__delay_1638___plus_1250;
  reg signed [16-1:0] __delay_data_1661__delay_1660__delay_1659___cond_1083;
  reg signed [16-1:0] __delay_data_1681__delay_1680__delay_1679___cond_1095;
  reg [16-1:0] __delay_data_1701__delay_1700__delay_1699___plus_1204;
  wire signed [64-1:0] __substreamoutput_data_1197;
  assign __substreamoutput_data_1197 = add_tree_3_sum_data;
  assign _acc_0_is_root = ((_stream_matmul_33_busy)? 0 : 1) && (((_stream_matmul_23_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1));
  assign _acc_0_stream_oready = ((_stream_matmul_33_busy)? _stream_matmul_33_stream_oready : 1) && (((_stream_matmul_23_busy)? _stream_matmul_23_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _acc_0_stream_internal_oready));
  wire signed [64-1:0] __substreamoutput_data_1218;
  assign __substreamoutput_data_1218 = add_tree_4_sum_data;
  reg [1-1:0] __variable_wdata_37;
  assign acc_1__reduce_reset_data = __variable_wdata_37;
  reg signed [64-1:0] __variable_wdata_22;
  assign acc_1_x_data = __variable_wdata_22;
  reg [7-1:0] __variable_wdata_23;
  assign acc_1_rshift_data = __variable_wdata_23;
  reg [32-1:0] __variable_wdata_24;
  assign acc_1_size_data = __variable_wdata_24;
  assign _acc_1_is_root = ((_stream_matmul_33_busy)? 0 : 1) && 1;
  assign _acc_1_stream_oready = ((_stream_matmul_33_busy)? _stream_matmul_33_stream_oready : 1) && _acc_1_stream_internal_oready;
  reg signed [16-1:0] __delay_data_1601__delay_1600__delay_1599___cond_1084;
  reg signed [16-1:0] __delay_data_1621__delay_1620__delay_1619___cond_1096;
  reg [16-1:0] __delay_data_1641__delay_1640__delay_1639___plus_1250;
  reg signed [16-1:0] __delay_data_1662__delay_1661__delay_1660___cond_1083;
  reg signed [16-1:0] __delay_data_1682__delay_1681__delay_1680___cond_1095;
  reg [16-1:0] __delay_data_1702__delay_1701__delay_1700___plus_1204;
  reg signed [16-1:0] __delay_data_1602__delay_1601__delay_1600___cond_1084;
  reg signed [16-1:0] __delay_data_1622__delay_1621__delay_1620___cond_1096;
  reg [16-1:0] __delay_data_1642__delay_1641__delay_1640___plus_1250;
  reg signed [16-1:0] __delay_data_1663__delay_1662__delay_1661___cond_1083;
  reg signed [16-1:0] __delay_data_1683__delay_1682__delay_1681___cond_1095;
  reg [16-1:0] __delay_data_1703__delay_1702__delay_1701___plus_1204;
  reg signed [16-1:0] __delay_data_1603__delay_1602__delay_1601___cond_1084;
  reg signed [16-1:0] __delay_data_1623__delay_1622__delay_1621___cond_1096;
  reg [16-1:0] __delay_data_1643__delay_1642__delay_1641___plus_1250;
  reg signed [16-1:0] __delay_data_1664__delay_1663__delay_1662___cond_1083;
  reg signed [16-1:0] __delay_data_1684__delay_1683__delay_1682___cond_1095;
  reg [16-1:0] __delay_data_1704__delay_1703__delay_1702___plus_1204;
  reg signed [16-1:0] __delay_data_1604__delay_1603__delay_1602___cond_1084;
  reg signed [16-1:0] __delay_data_1624__delay_1623__delay_1622___cond_1096;
  reg [16-1:0] __delay_data_1644__delay_1643__delay_1642___plus_1250;
  reg signed [16-1:0] __delay_data_1665__delay_1664__delay_1663___cond_1083;
  reg signed [16-1:0] __delay_data_1685__delay_1684__delay_1683___cond_1095;
  reg [16-1:0] __delay_data_1705__delay_1704__delay_1703___plus_1204;
  reg signed [16-1:0] __delay_data_1605__delay_1604__delay_1603___cond_1084;
  reg signed [16-1:0] __delay_data_1625__delay_1624__delay_1623___cond_1096;
  reg [16-1:0] __delay_data_1645__delay_1644__delay_1643___plus_1250;
  reg signed [16-1:0] __delay_data_1666__delay_1665__delay_1664___cond_1083;
  reg signed [16-1:0] __delay_data_1686__delay_1685__delay_1684___cond_1095;
  reg [16-1:0] __delay_data_1706__delay_1705__delay_1704___plus_1204;
  reg signed [16-1:0] __delay_data_1606__delay_1605__delay_1604___cond_1084;
  reg signed [16-1:0] __delay_data_1626__delay_1625__delay_1624___cond_1096;
  reg [16-1:0] __delay_data_1646__delay_1645__delay_1644___plus_1250;
  reg signed [16-1:0] __delay_data_1667__delay_1666__delay_1665___cond_1083;
  reg signed [16-1:0] __delay_data_1687__delay_1686__delay_1685___cond_1095;
  reg [16-1:0] __delay_data_1707__delay_1706__delay_1705___plus_1204;
  wire signed [64-1:0] __substreamoutput_data_1200;
  assign __substreamoutput_data_1200 = acc_0_sum_data;
  wire [1-1:0] __substreamoutput_data_1201;
  assign __substreamoutput_data_1201 = acc_0_valid_data;
  reg signed [64-1:0] _plus_data_1202;
  wire signed [64-1:0] __substreamoutput_data_1232;
  assign __substreamoutput_data_1232 = acc_1_sum_data;
  reg signed [64-1:0] _plus_data_1234;
  reg signed [16-1:0] __delay_data_1627__delay_1626__delay_1625___cond_1096;
  reg [16-1:0] __delay_data_1647__delay_1646__delay_1645___plus_1250;
  reg signed [16-1:0] __delay_data_1688__delay_1687__delay_1686___cond_1095;
  reg [16-1:0] __delay_data_1708__delay_1707__delay_1706___plus_1204;
  reg [1-1:0] __delay_data_1709__substreamoutput_1201;
  assign _mul_rshift_round_clip_6_is_root = ((_stream_matmul_33_busy)? 0 : 1) && (((_stream_matmul_23_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1));
  assign _mul_rshift_round_clip_6_stream_oready = ((_stream_matmul_33_busy)? _stream_matmul_33_stream_oready : 1) && (((_stream_matmul_23_busy)? _stream_matmul_23_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_rshift_round_clip_6_stream_internal_oready));
  reg signed [64-1:0] __variable_wdata_102;
  assign mul_rshift_round_clip_7_x_data = __variable_wdata_102;
  reg signed [16-1:0] __variable_wdata_103;
  assign mul_rshift_round_clip_7_y_data = __variable_wdata_103;
  reg [7-1:0] __variable_wdata_104;
  assign mul_rshift_round_clip_7_rshift_data = __variable_wdata_104;
  assign _mul_rshift_round_clip_7_is_root = ((_stream_matmul_33_busy)? 0 : 1) && 1;
  assign _mul_rshift_round_clip_7_stream_oready = ((_stream_matmul_33_busy)? _stream_matmul_33_stream_oready : 1) && _mul_rshift_round_clip_7_stream_internal_oready;
  assign _stream_matmul_33_stream_internal_oready = ((_stream_matmul_33_busy)? _mul_rshift_round_clip_7_stream_internal_oready : 1) && (((_stream_matmul_33_busy)? _mul_rshift_round_clip_6_stream_internal_oready : 1) && (((_stream_matmul_33_busy)? _acc_1_stream_internal_oready : 1) && (((_stream_matmul_33_busy)? _acc_0_stream_internal_oready : 1) && (((_stream_matmul_33_busy)? _add_tree_4_stream_internal_oready : 1) && (((_stream_matmul_33_busy)? _add_tree_3_stream_internal_oready : 1) && (((_stream_matmul_33_busy)? _mul_11_stream_internal_oready : 1) && (((_stream_matmul_33_busy)? _mul_10_stream_internal_oready : 1) && (((_stream_matmul_33_busy)? _mul_9_stream_internal_oready : 1) && (((_stream_matmul_33_busy)? _mul_8_stream_internal_oready : 1) && 1)))))))));
  reg [1-1:0] __delay_data_1710__delay_1709__substreamoutput_1201;
  reg [1-1:0] __delay_data_1711__delay_1710____substreamoutput_1201;
  reg [1-1:0] __delay_data_1712__delay_1711____substreamoutput_1201;
  reg [1-1:0] __delay_data_1713__delay_1712____substreamoutput_1201;
  reg [1-1:0] __delay_data_1714__delay_1713____substreamoutput_1201;
  reg [1-1:0] __delay_data_1715__delay_1714____substreamoutput_1201;
  reg [1-1:0] __delay_data_1716__delay_1715____substreamoutput_1201;
  reg [1-1:0] __delay_data_1717__delay_1716____substreamoutput_1201;
  reg [1-1:0] __delay_data_1718__delay_1717____substreamoutput_1201;
  wire signed [16-1:0] __substreamoutput_data_1205;
  assign __substreamoutput_data_1205 = mul_rshift_round_clip_6_z_data;
  wire signed [16-1:0] _reinterpretcast_src_1206;
  assign _reinterpretcast_src_1206 = __substreamoutput_data_1205;
  wire signed [16-1:0] _reinterpretcast_data_1206;
  assign _reinterpretcast_data_1206 = _reinterpretcast_src_1206;
  wire signed [16-1:0] __substreamoutput_data_1251;
  assign __substreamoutput_data_1251 = mul_rshift_round_clip_7_z_data;
  wire signed [16-1:0] _reinterpretcast_src_1252;
  assign _reinterpretcast_src_1252 = __substreamoutput_data_1251;
  wire signed [16-1:0] _reinterpretcast_data_1252;
  assign _reinterpretcast_data_1252 = _reinterpretcast_src_1252;
  wire [32-1:0] _cat_data_1253;
  assign _cat_data_1253 = { _reinterpretcast_data_1252, _reinterpretcast_data_1206 };
  wire [32-1:0] stream_matmul_33_sink_33_data;
  assign stream_matmul_33_sink_33_data = _cat_data_1253;
  wire [1-1:0] stream_matmul_33_sink_34_data;
  assign stream_matmul_33_sink_34_data = __delay_data_1718__delay_1717____substreamoutput_1201;
  wire _set_flag_1670;
  assign _set_flag_1670 = matmul_33_comp_fsm == 3;
  reg [9-1:0] __variable_wdata_1052;
  assign stream_matmul_33_parameter_0_data = __variable_wdata_1052;
  wire _set_flag_1671;
  assign _set_flag_1671 = matmul_33_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1053;
  assign stream_matmul_33_parameter_1_data = __variable_wdata_1053;
  wire _set_flag_1672;
  assign _set_flag_1672 = matmul_33_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1054;
  assign stream_matmul_33_parameter_2_data = __variable_wdata_1054;
  wire _set_flag_1673;
  assign _set_flag_1673 = matmul_33_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1055;
  assign stream_matmul_33_parameter_3_data = __variable_wdata_1055;
  wire _set_flag_1674;
  assign _set_flag_1674 = matmul_33_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_1056;
  assign stream_matmul_33_parameter_4_data = __variable_wdata_1056;
  wire _set_flag_1675;
  assign _set_flag_1675 = matmul_33_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1073;
  assign stream_matmul_33_parameter_6_data = __variable_wdata_1073;
  reg [32-1:0] _source_stream_matmul_33_source_7_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_33_source_7_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_33_source_7_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_33_source_7_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_33_source_7_pat_size_0;
  reg [33-1:0] _source_stream_matmul_33_source_7_pat_size_1;
  reg [33-1:0] _source_stream_matmul_33_source_7_pat_size_2;
  reg [33-1:0] _source_stream_matmul_33_source_7_pat_size_3;
  reg [32-1:0] _source_stream_matmul_33_source_7_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_33_source_7_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_33_source_7_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_33_source_7_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_33_source_7_pat_count_0;
  reg [33-1:0] _source_stream_matmul_33_source_7_pat_count_1;
  reg [33-1:0] _source_stream_matmul_33_source_7_pat_count_2;
  reg [33-1:0] _source_stream_matmul_33_source_7_pat_count_3;
  reg [33-1:0] _source_stream_matmul_33_source_7_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_33_source_7_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_33_source_7_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_33_source_7_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_33_source_7_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_33_source_7_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_33_source_7_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_33_source_7_pat_stride_buf_3;
  wire _set_flag_1676;
  assign _set_flag_1676 = matmul_33_comp_fsm == 3;
  assign ram_w32_l128_id1_0_addr = (_stream_matmul_33_stream_oready && _stream_matmul_33_source_7_source_ram_renable && (_stream_matmul_33_source_7_source_sel == 1))? _stream_matmul_33_source_7_source_ram_raddr : 'hx;
  assign ram_w32_l128_id1_0_enable = (_stream_matmul_33_stream_oready && _stream_matmul_33_source_7_source_ram_renable && (_stream_matmul_33_source_7_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_1677 = 1;
  wire [_tmp_1677-1:0] _tmp_1678;
  assign _tmp_1678 = _stream_matmul_33_stream_oready && _stream_matmul_33_source_7_source_ram_renable && (_stream_matmul_33_source_7_source_sel == 1);
  reg [_tmp_1677-1:0] __tmp_1678_1;
  assign _stream_matmul_33_source_7_source_ram_rdata = (_stream_matmul_33_source_7_source_sel == 1)? ram_w32_l128_id1_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1074;
  assign stream_matmul_33_source_7_data = __variable_wdata_1074;
  reg [32-1:0] _stream_matmul_33_source_7_source_pat_fsm_0;
  localparam _stream_matmul_33_source_7_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_matmul_33_source_7_source_pat_all_offset;
  assign _stream_matmul_33_source_7_source_pat_all_offset = _stream_matmul_33_source_7_source_offset_buf + _source_stream_matmul_33_source_7_pat_cur_offset_0 + _source_stream_matmul_33_source_7_pat_cur_offset_1 + _source_stream_matmul_33_source_7_pat_cur_offset_2 + _source_stream_matmul_33_source_7_pat_cur_offset_3;
  wire _set_flag_1679;
  assign _set_flag_1679 = matmul_33_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1085;
  assign stream_matmul_33_parameter_8_data = __variable_wdata_1085;
  reg [32-1:0] _source_stream_matmul_33_source_9_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_33_source_9_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_33_source_9_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_33_source_9_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_33_source_9_pat_size_0;
  reg [33-1:0] _source_stream_matmul_33_source_9_pat_size_1;
  reg [33-1:0] _source_stream_matmul_33_source_9_pat_size_2;
  reg [33-1:0] _source_stream_matmul_33_source_9_pat_size_3;
  reg [32-1:0] _source_stream_matmul_33_source_9_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_33_source_9_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_33_source_9_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_33_source_9_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_33_source_9_pat_count_0;
  reg [33-1:0] _source_stream_matmul_33_source_9_pat_count_1;
  reg [33-1:0] _source_stream_matmul_33_source_9_pat_count_2;
  reg [33-1:0] _source_stream_matmul_33_source_9_pat_count_3;
  reg [33-1:0] _source_stream_matmul_33_source_9_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_33_source_9_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_33_source_9_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_33_source_9_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_33_source_9_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_33_source_9_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_33_source_9_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_33_source_9_pat_stride_buf_3;
  wire _set_flag_1680;
  assign _set_flag_1680 = matmul_33_comp_fsm == 3;
  assign ram_w32_l128_id2_0_addr = (_stream_matmul_33_stream_oready && _stream_matmul_33_source_9_source_ram_renable && (_stream_matmul_33_source_9_source_sel == 2))? _stream_matmul_33_source_9_source_ram_raddr : 'hx;
  assign ram_w32_l128_id2_0_enable = (_stream_matmul_33_stream_oready && _stream_matmul_33_source_9_source_ram_renable && (_stream_matmul_33_source_9_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_1681 = 1;
  wire [_tmp_1681-1:0] _tmp_1682;
  assign _tmp_1682 = _stream_matmul_33_stream_oready && _stream_matmul_33_source_9_source_ram_renable && (_stream_matmul_33_source_9_source_sel == 2);
  reg [_tmp_1681-1:0] __tmp_1682_1;
  assign _stream_matmul_33_source_9_source_ram_rdata = (_stream_matmul_33_source_9_source_sel == 2)? ram_w32_l128_id2_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1086;
  assign stream_matmul_33_source_9_data = __variable_wdata_1086;
  reg [32-1:0] _stream_matmul_33_source_9_source_pat_fsm_1;
  localparam _stream_matmul_33_source_9_source_pat_fsm_1_init = 0;
  wire [32-1:0] _stream_matmul_33_source_9_source_pat_all_offset;
  assign _stream_matmul_33_source_9_source_pat_all_offset = _stream_matmul_33_source_9_source_offset_buf + _source_stream_matmul_33_source_9_pat_cur_offset_0 + _source_stream_matmul_33_source_9_pat_cur_offset_1 + _source_stream_matmul_33_source_9_pat_cur_offset_2 + _source_stream_matmul_33_source_9_pat_cur_offset_3;
  wire _set_flag_1683;
  assign _set_flag_1683 = matmul_33_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1097;
  assign stream_matmul_33_parameter_10_data = __variable_wdata_1097;
  wire _set_flag_1684;
  assign _set_flag_1684 = matmul_33_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_1098;
  assign stream_matmul_33_source_11_data = __variable_wdata_1098;
  wire _set_flag_1685;
  assign _set_flag_1685 = matmul_33_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1109;
  assign stream_matmul_33_parameter_12_data = __variable_wdata_1109;
  wire _set_flag_1686;
  assign _set_flag_1686 = matmul_33_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_1110;
  assign stream_matmul_33_source_13_data = __variable_wdata_1110;
  wire _set_flag_1687;
  assign _set_flag_1687 = matmul_33_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1121;
  assign stream_matmul_33_parameter_14_data = __variable_wdata_1121;
  wire _set_flag_1688;
  assign _set_flag_1688 = matmul_33_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_1122;
  assign stream_matmul_33_source_15_data = __variable_wdata_1122;
  wire _set_flag_1689;
  assign _set_flag_1689 = matmul_33_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1133;
  assign stream_matmul_33_parameter_16_data = __variable_wdata_1133;
  wire _set_flag_1690;
  assign _set_flag_1690 = matmul_33_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1134;
  assign stream_matmul_33_parameter_17_data = __variable_wdata_1134;
  wire _set_flag_1691;
  assign _set_flag_1691 = matmul_33_comp_fsm == 3;
  reg [5-1:0] __variable_wdata_1135;
  assign stream_matmul_33_parameter_18_data = __variable_wdata_1135;
  wire _set_flag_1692;
  assign _set_flag_1692 = matmul_33_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1136;
  assign stream_matmul_33_parameter_19_data = __variable_wdata_1136;
  reg [32-1:0] _source_stream_matmul_33_source_20_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_33_source_20_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_33_source_20_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_33_source_20_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_33_source_20_pat_size_0;
  reg [33-1:0] _source_stream_matmul_33_source_20_pat_size_1;
  reg [33-1:0] _source_stream_matmul_33_source_20_pat_size_2;
  reg [33-1:0] _source_stream_matmul_33_source_20_pat_size_3;
  reg [32-1:0] _source_stream_matmul_33_source_20_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_33_source_20_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_33_source_20_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_33_source_20_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_33_source_20_pat_count_0;
  reg [33-1:0] _source_stream_matmul_33_source_20_pat_count_1;
  reg [33-1:0] _source_stream_matmul_33_source_20_pat_count_2;
  reg [33-1:0] _source_stream_matmul_33_source_20_pat_count_3;
  reg [33-1:0] _source_stream_matmul_33_source_20_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_33_source_20_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_33_source_20_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_33_source_20_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_33_source_20_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_33_source_20_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_33_source_20_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_33_source_20_pat_stride_buf_3;
  wire _set_flag_1693;
  assign _set_flag_1693 = matmul_33_comp_fsm == 3;
  assign ram_w32_l512_id0_0_addr = (_stream_matmul_33_stream_oready && _stream_matmul_33_source_20_source_ram_renable && (_stream_matmul_33_source_20_source_sel == 3))? _stream_matmul_33_source_20_source_ram_raddr : 'hx;
  assign ram_w32_l512_id0_0_enable = (_stream_matmul_33_stream_oready && _stream_matmul_33_source_20_source_ram_renable && (_stream_matmul_33_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1694 = 1;
  wire [_tmp_1694-1:0] _tmp_1695;
  assign _tmp_1695 = _stream_matmul_33_stream_oready && _stream_matmul_33_source_20_source_ram_renable && (_stream_matmul_33_source_20_source_sel == 3);
  reg [_tmp_1694-1:0] __tmp_1695_1;
  assign _stream_matmul_33_source_20_source_ram_rdata = (_stream_matmul_33_source_20_source_sel == 3)? ram_w32_l512_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1137;
  assign stream_matmul_33_source_20_data = __variable_wdata_1137;
  reg [32-1:0] _stream_matmul_33_source_20_source_pat_fsm_2;
  localparam _stream_matmul_33_source_20_source_pat_fsm_2_init = 0;
  wire [32-1:0] _stream_matmul_33_source_20_source_pat_all_offset;
  assign _stream_matmul_33_source_20_source_pat_all_offset = _stream_matmul_33_source_20_source_offset_buf + _source_stream_matmul_33_source_20_pat_cur_offset_0 + _source_stream_matmul_33_source_20_pat_cur_offset_1 + _source_stream_matmul_33_source_20_pat_cur_offset_2 + _source_stream_matmul_33_source_20_pat_cur_offset_3;
  reg [32-1:0] _source_stream_matmul_33_source_21_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_33_source_21_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_33_source_21_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_33_source_21_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_33_source_21_pat_size_0;
  reg [33-1:0] _source_stream_matmul_33_source_21_pat_size_1;
  reg [33-1:0] _source_stream_matmul_33_source_21_pat_size_2;
  reg [33-1:0] _source_stream_matmul_33_source_21_pat_size_3;
  reg [32-1:0] _source_stream_matmul_33_source_21_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_33_source_21_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_33_source_21_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_33_source_21_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_33_source_21_pat_count_0;
  reg [33-1:0] _source_stream_matmul_33_source_21_pat_count_1;
  reg [33-1:0] _source_stream_matmul_33_source_21_pat_count_2;
  reg [33-1:0] _source_stream_matmul_33_source_21_pat_count_3;
  reg [33-1:0] _source_stream_matmul_33_source_21_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_33_source_21_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_33_source_21_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_33_source_21_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_33_source_21_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_33_source_21_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_33_source_21_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_33_source_21_pat_stride_buf_3;
  wire _set_flag_1696;
  assign _set_flag_1696 = matmul_33_comp_fsm == 3;
  assign ram_w32_l512_id1_0_addr = (_stream_matmul_33_stream_oready && _stream_matmul_33_source_21_source_ram_renable && (_stream_matmul_33_source_21_source_sel == 4))? _stream_matmul_33_source_21_source_ram_raddr : 'hx;
  assign ram_w32_l512_id1_0_enable = (_stream_matmul_33_stream_oready && _stream_matmul_33_source_21_source_ram_renable && (_stream_matmul_33_source_21_source_sel == 4))? 1'd1 : 0;
  localparam _tmp_1697 = 1;
  wire [_tmp_1697-1:0] _tmp_1698;
  assign _tmp_1698 = _stream_matmul_33_stream_oready && _stream_matmul_33_source_21_source_ram_renable && (_stream_matmul_33_source_21_source_sel == 4);
  reg [_tmp_1697-1:0] __tmp_1698_1;
  assign _stream_matmul_33_source_21_source_ram_rdata = (_stream_matmul_33_source_21_source_sel == 4)? ram_w32_l512_id1_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1158;
  assign stream_matmul_33_source_21_data = __variable_wdata_1158;
  reg [32-1:0] _stream_matmul_33_source_21_source_pat_fsm_3;
  localparam _stream_matmul_33_source_21_source_pat_fsm_3_init = 0;
  wire [32-1:0] _stream_matmul_33_source_21_source_pat_all_offset;
  assign _stream_matmul_33_source_21_source_pat_all_offset = _stream_matmul_33_source_21_source_offset_buf + _source_stream_matmul_33_source_21_pat_cur_offset_0 + _source_stream_matmul_33_source_21_pat_cur_offset_1 + _source_stream_matmul_33_source_21_pat_cur_offset_2 + _source_stream_matmul_33_source_21_pat_cur_offset_3;
  reg [32-1:0] _source_stream_matmul_33_source_22_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_33_source_22_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_33_source_22_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_33_source_22_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_33_source_22_pat_size_0;
  reg [33-1:0] _source_stream_matmul_33_source_22_pat_size_1;
  reg [33-1:0] _source_stream_matmul_33_source_22_pat_size_2;
  reg [33-1:0] _source_stream_matmul_33_source_22_pat_size_3;
  reg [32-1:0] _source_stream_matmul_33_source_22_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_33_source_22_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_33_source_22_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_33_source_22_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_33_source_22_pat_count_0;
  reg [33-1:0] _source_stream_matmul_33_source_22_pat_count_1;
  reg [33-1:0] _source_stream_matmul_33_source_22_pat_count_2;
  reg [33-1:0] _source_stream_matmul_33_source_22_pat_count_3;
  reg [33-1:0] _source_stream_matmul_33_source_22_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_33_source_22_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_33_source_22_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_33_source_22_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_33_source_22_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_33_source_22_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_33_source_22_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_33_source_22_pat_stride_buf_3;
  wire _set_flag_1699;
  assign _set_flag_1699 = matmul_33_comp_fsm == 3;
  assign ram_w32_l1024_id0_0_addr = (_stream_matmul_33_stream_oready && _stream_matmul_33_source_22_source_ram_renable && (_stream_matmul_33_source_22_source_sel == 5))? _stream_matmul_33_source_22_source_ram_raddr : 
                                    (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_6_sink_wenable && (_stream_max_pool_serial_6_sink_6_sink_sel == 2))? _stream_max_pool_serial_6_sink_6_sink_waddr : 'hx;
  assign ram_w32_l1024_id0_0_enable = (_stream_matmul_33_stream_oready && _stream_matmul_33_source_22_source_ram_renable && (_stream_matmul_33_source_22_source_sel == 5))? 1'd1 : 
                                      (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_6_sink_wenable && (_stream_max_pool_serial_6_sink_6_sink_sel == 2))? 1'd1 : 0;
  localparam _tmp_1700 = 1;
  wire [_tmp_1700-1:0] _tmp_1701;
  assign _tmp_1701 = _stream_matmul_33_stream_oready && _stream_matmul_33_source_22_source_ram_renable && (_stream_matmul_33_source_22_source_sel == 5);
  reg [_tmp_1700-1:0] __tmp_1701_1;
  assign _stream_matmul_33_source_22_source_ram_rdata = (_stream_matmul_33_source_22_source_sel == 5)? ram_w32_l1024_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1159;
  assign stream_matmul_33_source_22_data = __variable_wdata_1159;
  reg [32-1:0] _stream_matmul_33_source_22_source_pat_fsm_4;
  localparam _stream_matmul_33_source_22_source_pat_fsm_4_init = 0;
  wire [32-1:0] _stream_matmul_33_source_22_source_pat_all_offset;
  assign _stream_matmul_33_source_22_source_pat_all_offset = _stream_matmul_33_source_22_source_offset_buf + _source_stream_matmul_33_source_22_pat_cur_offset_0 + _source_stream_matmul_33_source_22_pat_cur_offset_1 + _source_stream_matmul_33_source_22_pat_cur_offset_2 + _source_stream_matmul_33_source_22_pat_cur_offset_3;
  wire _set_flag_1702;
  assign _set_flag_1702 = matmul_33_comp_fsm == 3;
  reg _tmp_1703;
  reg _tmp_1704;
  reg _tmp_1705;
  reg _tmp_1706;
  reg _tmp_1707;
  reg _tmp_1708;
  reg _tmp_1709;
  reg _tmp_1710;
  reg _tmp_1711;
  reg _tmp_1712;
  reg _tmp_1713;
  reg _tmp_1714;
  reg _tmp_1715;
  reg _tmp_1716;
  reg _tmp_1717;
  reg _tmp_1718;
  reg _tmp_1719;
  reg _tmp_1720;
  reg _tmp_1721;
  reg _tmp_1722;
  reg _tmp_1723;
  reg _tmp_1724;
  reg _tmp_1725;
  reg _tmp_1726;
  reg _tmp_1727;
  reg _tmp_1728;
  reg _tmp_1729;
  reg _tmp_1730;
  reg _tmp_1731;
  reg _tmp_1732;
  reg _tmp_1733;
  reg _tmp_1734;
  localparam _tmp_1735 = 33;
  wire [_tmp_1735-1:0] _tmp_1736;
  assign _tmp_1736 = matmul_33_stream_out_local + matmul_33_out_page_comp_offset_buf;
  reg [_tmp_1735-1:0] _tmp_1737;
  reg [_tmp_1735-1:0] _tmp_1738;
  reg [_tmp_1735-1:0] _tmp_1739;
  reg [_tmp_1735-1:0] _tmp_1740;
  reg [_tmp_1735-1:0] _tmp_1741;
  reg [_tmp_1735-1:0] _tmp_1742;
  reg [_tmp_1735-1:0] _tmp_1743;
  reg [_tmp_1735-1:0] _tmp_1744;
  reg [_tmp_1735-1:0] _tmp_1745;
  reg [_tmp_1735-1:0] _tmp_1746;
  reg [_tmp_1735-1:0] _tmp_1747;
  reg [_tmp_1735-1:0] _tmp_1748;
  reg [_tmp_1735-1:0] _tmp_1749;
  reg [_tmp_1735-1:0] _tmp_1750;
  reg [_tmp_1735-1:0] _tmp_1751;
  reg [_tmp_1735-1:0] _tmp_1752;
  reg [_tmp_1735-1:0] _tmp_1753;
  reg [_tmp_1735-1:0] _tmp_1754;
  reg [_tmp_1735-1:0] _tmp_1755;
  reg [_tmp_1735-1:0] _tmp_1756;
  reg [_tmp_1735-1:0] _tmp_1757;
  reg [_tmp_1735-1:0] _tmp_1758;
  reg [_tmp_1735-1:0] _tmp_1759;
  reg [_tmp_1735-1:0] _tmp_1760;
  reg [_tmp_1735-1:0] _tmp_1761;
  reg [_tmp_1735-1:0] _tmp_1762;
  reg [_tmp_1735-1:0] _tmp_1763;
  reg [_tmp_1735-1:0] _tmp_1764;
  reg [_tmp_1735-1:0] _tmp_1765;
  reg [_tmp_1735-1:0] _tmp_1766;
  reg [_tmp_1735-1:0] _tmp_1767;
  reg [_tmp_1735-1:0] _tmp_1768;
  reg [32-1:0] _tmp_1769;
  reg [32-1:0] _tmp_1770;
  reg [32-1:0] _tmp_1771;
  reg [32-1:0] _tmp_1772;
  reg [32-1:0] _tmp_1773;
  reg [32-1:0] _tmp_1774;
  reg [32-1:0] _tmp_1775;
  reg [32-1:0] _tmp_1776;
  reg [32-1:0] _tmp_1777;
  reg [32-1:0] _tmp_1778;
  reg [32-1:0] _tmp_1779;
  reg [32-1:0] _tmp_1780;
  reg [32-1:0] _tmp_1781;
  reg [32-1:0] _tmp_1782;
  reg [32-1:0] _tmp_1783;
  reg [32-1:0] _tmp_1784;
  reg [32-1:0] _tmp_1785;
  reg [32-1:0] _tmp_1786;
  reg [32-1:0] _tmp_1787;
  reg [32-1:0] _tmp_1788;
  reg [32-1:0] _tmp_1789;
  reg [32-1:0] _tmp_1790;
  reg [32-1:0] _tmp_1791;
  reg [32-1:0] _tmp_1792;
  reg [32-1:0] _tmp_1793;
  reg [32-1:0] _tmp_1794;
  reg [32-1:0] _tmp_1795;
  reg [32-1:0] _tmp_1796;
  reg [32-1:0] _tmp_1797;
  reg [32-1:0] _tmp_1798;
  reg [32-1:0] _tmp_1799;
  reg [32-1:0] _tmp_1800;
  assign ram_w32_l128_id0_0_addr = (_stream_matmul_33_stream_oready && _stream_matmul_33_sink_33_sink_wenable && (_stream_matmul_33_sink_33_sink_sel == 6))? _stream_matmul_33_sink_33_sink_waddr : 'hx;
  assign ram_w32_l128_id0_0_wdata = (_stream_matmul_33_stream_oready && _stream_matmul_33_sink_33_sink_wenable && (_stream_matmul_33_sink_33_sink_sel == 6))? _stream_matmul_33_sink_33_sink_wdata : 'hx;
  assign ram_w32_l128_id0_0_wenable = (_stream_matmul_33_stream_oready && _stream_matmul_33_sink_33_sink_wenable && (_stream_matmul_33_sink_33_sink_sel == 6))? 1'd1 : 0;
  assign ram_w32_l128_id0_0_enable = (_stream_matmul_33_stream_oready && _stream_matmul_33_sink_33_sink_wenable && (_stream_matmul_33_sink_33_sink_sel == 6))? 1'd1 : 0;
  reg [32-1:0] _stream_matmul_33_sink_33_sink_fsm_5;
  localparam _stream_matmul_33_sink_33_sink_fsm_5_init = 0;
  wire _set_flag_1801;
  assign _set_flag_1801 = matmul_33_comp_fsm == 4;
  assign _stream_matmul_33_run_flag = (_set_flag_1801)? 1 : 0;
  reg _tmp_1802;
  reg _tmp_1803;
  reg _tmp_1804;
  assign _add_tree_3_source_stop = _add_tree_3_stream_oready && 1'd0;
  reg _tmp_1805;
  reg _tmp_1806;
  reg _tmp_1807;
  assign _add_tree_3_sink_start = _tmp_1807;
  reg _tmp_1808;
  reg _tmp_1809;
  reg _tmp_1810;
  assign _add_tree_3_sink_stop = _tmp_1810;
  reg _tmp_1811;
  reg _tmp_1812;
  reg _tmp_1813;
  assign _add_tree_3_sink_busy = _tmp_1813;
  reg _tmp_1814;
  assign _add_tree_3_busy = _add_tree_3_source_busy || _add_tree_3_sink_busy || _add_tree_3_busy_reg;
  reg _tmp_1815;
  reg _tmp_1816;
  reg _tmp_1817;
  assign _add_tree_4_source_stop = _add_tree_4_stream_oready && 1'd0;
  reg _tmp_1818;
  reg _tmp_1819;
  reg _tmp_1820;
  assign _add_tree_4_sink_start = _tmp_1820;
  reg _tmp_1821;
  reg _tmp_1822;
  reg _tmp_1823;
  assign _add_tree_4_sink_stop = _tmp_1823;
  reg _tmp_1824;
  reg _tmp_1825;
  reg _tmp_1826;
  assign _add_tree_4_sink_busy = _tmp_1826;
  reg _tmp_1827;
  assign _add_tree_4_busy = _add_tree_4_source_busy || _add_tree_4_sink_busy || _add_tree_4_busy_reg;
  reg _tmp_1828;
  reg _tmp_1829;
  reg _tmp_1830;
  reg _tmp_1831;
  reg _tmp_1832;
  reg _tmp_1833;
  reg _tmp_1834;
  reg _tmp_1835;
  reg _tmp_1836;
  reg _tmp_1837;
  assign _acc_1_source_stop = _acc_1_stream_oready && 1'd0;
  reg _tmp_1838;
  reg _tmp_1839;
  reg _tmp_1840;
  reg _tmp_1841;
  reg _tmp_1842;
  reg _tmp_1843;
  reg _tmp_1844;
  assign _acc_1_sink_start = _tmp_1844;
  reg _tmp_1845;
  reg _tmp_1846;
  reg _tmp_1847;
  reg _tmp_1848;
  reg _tmp_1849;
  reg _tmp_1850;
  reg _tmp_1851;
  assign _acc_1_sink_stop = _tmp_1851;
  reg _tmp_1852;
  reg _tmp_1853;
  reg _tmp_1854;
  reg _tmp_1855;
  reg _tmp_1856;
  reg _tmp_1857;
  reg _tmp_1858;
  assign _acc_1_sink_busy = _tmp_1858;
  reg _tmp_1859;
  assign _acc_1_busy = _acc_1_source_busy || _acc_1_sink_busy || _acc_1_busy_reg;
  reg _tmp_1860;
  reg _tmp_1861;
  reg _tmp_1862;
  assign _mul_rshift_round_clip_7_source_stop = _mul_rshift_round_clip_7_stream_oready && 1'd0;
  reg _tmp_1863;
  reg _tmp_1864;
  reg _tmp_1865;
  reg _tmp_1866;
  reg _tmp_1867;
  reg _tmp_1868;
  reg _tmp_1869;
  reg _tmp_1870;
  reg _tmp_1871;
  reg _tmp_1872;
  assign _mul_rshift_round_clip_7_sink_start = _tmp_1872;
  reg _tmp_1873;
  reg _tmp_1874;
  reg _tmp_1875;
  reg _tmp_1876;
  reg _tmp_1877;
  reg _tmp_1878;
  reg _tmp_1879;
  reg _tmp_1880;
  reg _tmp_1881;
  reg _tmp_1882;
  assign _mul_rshift_round_clip_7_sink_stop = _tmp_1882;
  reg _tmp_1883;
  reg _tmp_1884;
  reg _tmp_1885;
  reg _tmp_1886;
  reg _tmp_1887;
  reg _tmp_1888;
  reg _tmp_1889;
  reg _tmp_1890;
  reg _tmp_1891;
  reg _tmp_1892;
  assign _mul_rshift_round_clip_7_sink_busy = _tmp_1892;
  reg _tmp_1893;
  assign _mul_rshift_round_clip_7_busy = _mul_rshift_round_clip_7_source_busy || _mul_rshift_round_clip_7_sink_busy || _mul_rshift_round_clip_7_busy_reg;
  reg _tmp_1894;
  reg _tmp_1895;
  reg _tmp_1896;
  reg _tmp_1897;
  reg _tmp_1898;
  reg _tmp_1899;
  reg [1-1:0] __variable_wdata_1057;
  assign stream_matmul_33__reduce_reset_data = __variable_wdata_1057;
  reg _tmp_1900;
  reg _tmp_1901;
  reg _tmp_1902;
  reg _tmp_1903;
  assign _stream_matmul_33_source_stop = _stream_matmul_33_stream_oready && (_stream_matmul_33_source_11_idle && _stream_matmul_33_source_13_idle && _stream_matmul_33_source_15_idle && _stream_matmul_33_source_20_idle && _stream_matmul_33_source_21_idle && _stream_matmul_33_source_22_idle && _stream_matmul_33_source_7_idle && _stream_matmul_33_source_9_idle && (_stream_matmul_33_fsm == 3));
  localparam _tmp_1904 = 1;
  wire [_tmp_1904-1:0] _tmp_1905;
  assign _tmp_1905 = _stream_matmul_33_source_11_idle && _stream_matmul_33_source_13_idle && _stream_matmul_33_source_15_idle && _stream_matmul_33_source_20_idle && _stream_matmul_33_source_21_idle && _stream_matmul_33_source_22_idle && _stream_matmul_33_source_7_idle && _stream_matmul_33_source_9_idle && (_stream_matmul_33_fsm == 3);
  reg [_tmp_1904-1:0] _tmp_1906;
  localparam _tmp_1907 = 1;
  wire [_tmp_1907-1:0] _tmp_1908;
  assign _tmp_1908 = _stream_matmul_33_source_11_idle && _stream_matmul_33_source_13_idle && _stream_matmul_33_source_15_idle && _stream_matmul_33_source_20_idle && _stream_matmul_33_source_21_idle && _stream_matmul_33_source_22_idle && _stream_matmul_33_source_7_idle && _stream_matmul_33_source_9_idle && (_stream_matmul_33_fsm == 3);
  reg [_tmp_1907-1:0] _tmp_1909;
  reg _tmp_1910;
  reg _tmp_1911;
  reg _tmp_1912;
  reg _tmp_1913;
  reg _tmp_1914;
  reg _tmp_1915;
  reg _tmp_1916;
  reg _tmp_1917;
  reg _tmp_1918;
  reg _tmp_1919;
  reg _tmp_1920;
  reg _tmp_1921;
  reg _tmp_1922;
  reg _tmp_1923;
  reg _tmp_1924;
  reg _tmp_1925;
  reg _tmp_1926;
  reg _tmp_1927;
  reg _tmp_1928;
  reg _tmp_1929;
  reg _tmp_1930;
  reg _tmp_1931;
  reg _tmp_1932;
  reg _tmp_1933;
  reg _tmp_1934;
  reg _tmp_1935;
  reg _tmp_1936;
  reg _tmp_1937;
  reg _tmp_1938;
  reg _tmp_1939;
  reg _tmp_1940;
  reg _tmp_1941;
  assign _stream_matmul_33_sink_start = _tmp_1941;
  reg _tmp_1942;
  reg _tmp_1943;
  reg _tmp_1944;
  reg _tmp_1945;
  reg _tmp_1946;
  reg _tmp_1947;
  reg _tmp_1948;
  reg _tmp_1949;
  reg _tmp_1950;
  reg _tmp_1951;
  reg _tmp_1952;
  reg _tmp_1953;
  reg _tmp_1954;
  reg _tmp_1955;
  reg _tmp_1956;
  reg _tmp_1957;
  reg _tmp_1958;
  reg _tmp_1959;
  reg _tmp_1960;
  reg _tmp_1961;
  reg _tmp_1962;
  reg _tmp_1963;
  reg _tmp_1964;
  reg _tmp_1965;
  reg _tmp_1966;
  reg _tmp_1967;
  reg _tmp_1968;
  reg _tmp_1969;
  reg _tmp_1970;
  reg _tmp_1971;
  reg _tmp_1972;
  reg _tmp_1973;
  assign _stream_matmul_33_sink_stop = _tmp_1973;
  reg _tmp_1974;
  reg _tmp_1975;
  reg _tmp_1976;
  reg _tmp_1977;
  reg _tmp_1978;
  reg _tmp_1979;
  reg _tmp_1980;
  reg _tmp_1981;
  reg _tmp_1982;
  reg _tmp_1983;
  reg _tmp_1984;
  reg _tmp_1985;
  reg _tmp_1986;
  reg _tmp_1987;
  reg _tmp_1988;
  reg _tmp_1989;
  reg _tmp_1990;
  reg _tmp_1991;
  reg _tmp_1992;
  reg _tmp_1993;
  reg _tmp_1994;
  reg _tmp_1995;
  reg _tmp_1996;
  reg _tmp_1997;
  reg _tmp_1998;
  reg _tmp_1999;
  reg _tmp_2000;
  reg _tmp_2001;
  reg _tmp_2002;
  reg _tmp_2003;
  reg _tmp_2004;
  reg _tmp_2005;
  assign _stream_matmul_33_sink_busy = _tmp_2005;
  reg _tmp_2006;
  assign _stream_matmul_33_busy = _stream_matmul_33_source_busy || _stream_matmul_33_sink_busy || _stream_matmul_33_busy_reg;
  wire matmul_33_dma_out_mask_0;
  assign matmul_33_dma_out_mask_0 = matmul_33_out_row_count + 0 >= cparam_matmul_33_out_num_row;
  wire [32-1:0] mask_addr_shifted_2007;
  assign mask_addr_shifted_2007 = matmul_33_objaddr + (matmul_33_out_base_offset + cparam_matmul_33_out_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_2008;
  assign mask_addr_masked_2008 = mask_addr_shifted_2007 << 2;
  reg [32-1:0] read_burst_fsm_37;
  localparam read_burst_fsm_37_init = 0;
  reg [7-1:0] read_burst_addr_2009;
  reg [7-1:0] read_burst_stride_2010;
  reg [33-1:0] read_burst_length_2011;
  reg read_burst_rvalid_2012;
  reg read_burst_rlast_2013;
  assign ram_w32_l128_id0_1_addr = ((read_burst_fsm_37 == 1) && (!read_burst_rvalid_2012 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_addr_2009 : 'hx;
  assign ram_w32_l128_id0_1_enable = ((read_burst_fsm_37 == 1) && (!read_burst_rvalid_2012 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  localparam _tmp_2014 = 1;
  wire [_tmp_2014-1:0] _tmp_2015;
  assign _tmp_2015 = (read_burst_fsm_37 == 1) && (!read_burst_rvalid_2012 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_2014-1:0] __tmp_2015_1;
  wire [32-1:0] read_burst_rdata_2016;
  assign read_burst_rdata_2016 = ram_w32_l128_id0_1_rdata;
  assign _maxi_write_req_fifo_deq = ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1)) && !_maxi_write_req_fifo_empty)? 1 : 0;
  reg _maxi_wdata_cond_2_1;
  wire matmul_33_update_filter;
  assign matmul_33_update_filter = (cparam_matmul_33_data_stationary == 0) && (matmul_33_row_count >= cparam_matmul_33_max_row_count) && (matmul_33_bat_count >= cparam_matmul_33_max_bat_count) || (cparam_matmul_33_data_stationary == 1) && !cparam_matmul_33_keep_filter;
  wire matmul_33_update_act;
  assign matmul_33_update_act = (cparam_matmul_33_data_stationary == 1) && (matmul_33_och_count >= cparam_matmul_33_max_och_count) || (cparam_matmul_33_data_stationary == 0);
  wire matmul_33_mux_next_dma_flag_0;
  assign matmul_33_mux_next_dma_flag_0 = (matmul_33_row_select == 0)? (matmul_33_row_count >= cparam_matmul_33_max_row_count)? 1 : cparam_matmul_33_dma_flag_conds_0 : 1'd0;

  always @(posedge CLK) begin
    _RESETN_inv_1 <= RESETN_inv;
    _RESETN_inv_2 <= _RESETN_inv_1;
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      maxi_awaddr <= 0;
      maxi_awlen <= 0;
      maxi_awvalid <= 0;
      _maxi_waddr_cond_0_1 <= 0;
    end else begin
      if(_maxi_waddr_cond_0_1) begin
        maxi_awvalid <= 0;
      end 
      if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (_maxi_outstanding_wcount < 6) && ((_maxi_outstanding_wcount < 6) && (maxi_awready || !maxi_awvalid))) begin
        maxi_awaddr <= _maxi_write_global_addr;
        maxi_awlen <= _maxi_write_cur_global_size - 1;
        maxi_awvalid <= 1;
      end 
      if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (_maxi_outstanding_wcount < 6) && ((_maxi_outstanding_wcount < 6) && (maxi_awready || !maxi_awvalid)) && (_maxi_write_cur_global_size == 0)) begin
        maxi_awvalid <= 0;
      end 
      _maxi_waddr_cond_0_1 <= 1;
      if(maxi_awvalid && !maxi_awready) begin
        maxi_awvalid <= maxi_awvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_wdata_sb_0 <= 0;
      _maxi_wvalid_sb_0 <= 0;
      _maxi_wlast_sb_0 <= 0;
      _maxi_wstrb_sb_0 <= 0;
      _maxi_wdata_cond_0_1 <= 0;
      _maxi_wdata_cond_1_1 <= 0;
      _maxi_wdata_cond_2_1 <= 0;
    end else begin
      if(_maxi_wdata_cond_0_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if(_maxi_wdata_cond_1_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if(_maxi_wdata_cond_2_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if((_maxi_write_op_sel_buf == 1) && read_burst_packed_rvalid_1169 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_packed_rdata_1179;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_packed_rlast_1170 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_0_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
      if((_maxi_write_op_sel_buf == 2) && read_burst_rvalid_1301 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_rdata_1305;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_rlast_1302 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_1_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
      if((_maxi_write_op_sel_buf == 3) && read_burst_rvalid_2012 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_rdata_2016;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_rlast_2013 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_2_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _sb_maxi_writedata_data_6 <= 0;
      _sb_maxi_writedata_valid_7 <= 0;
      _sb_maxi_writedata_tmp_data_9 <= 0;
      _sb_maxi_writedata_tmp_valid_10 <= 0;
    end else begin
      if(_sb_maxi_writedata_m_ready_5 || !_sb_maxi_writedata_valid_7) begin
        _sb_maxi_writedata_data_6 <= _sb_maxi_writedata_next_data_11;
        _sb_maxi_writedata_valid_7 <= _sb_maxi_writedata_next_valid_12;
      end 
      if(!_sb_maxi_writedata_tmp_valid_10 && _sb_maxi_writedata_valid_7 && !_sb_maxi_writedata_m_ready_5) begin
        _sb_maxi_writedata_tmp_data_9 <= _sb_maxi_writedata_s_data_3;
        _sb_maxi_writedata_tmp_valid_10 <= _sb_maxi_writedata_s_valid_4;
      end 
      if(_sb_maxi_writedata_tmp_valid_10 && _sb_maxi_writedata_m_ready_5) begin
        _sb_maxi_writedata_tmp_valid_10 <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      maxi_araddr <= 0;
      maxi_arlen <= 0;
      maxi_arvalid <= 0;
      _maxi_raddr_cond_0_1 <= 0;
    end else begin
      if(_maxi_raddr_cond_0_1) begin
        maxi_arvalid <= 0;
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid)) begin
        maxi_araddr <= _maxi_read_global_addr;
        maxi_arlen <= _maxi_read_cur_global_size - 1;
        maxi_arvalid <= 1;
      end 
      _maxi_raddr_cond_0_1 <= 1;
      if(maxi_arvalid && !maxi_arready) begin
        maxi_arvalid <= maxi_arvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _sb_maxi_readdata_data_21 <= 0;
      _sb_maxi_readdata_valid_22 <= 0;
      _sb_maxi_readdata_tmp_data_24 <= 0;
      _sb_maxi_readdata_tmp_valid_25 <= 0;
    end else begin
      if(_sb_maxi_readdata_m_ready_20 || !_sb_maxi_readdata_valid_22) begin
        _sb_maxi_readdata_data_21 <= _sb_maxi_readdata_next_data_26;
        _sb_maxi_readdata_valid_22 <= _sb_maxi_readdata_next_valid_27;
      end 
      if(!_sb_maxi_readdata_tmp_valid_25 && _sb_maxi_readdata_valid_22 && !_sb_maxi_readdata_m_ready_20) begin
        _sb_maxi_readdata_tmp_data_24 <= _sb_maxi_readdata_s_data_18;
        _sb_maxi_readdata_tmp_valid_25 <= _sb_maxi_readdata_s_valid_19;
      end 
      if(_sb_maxi_readdata_tmp_valid_25 && _sb_maxi_readdata_m_ready_20) begin
        _sb_maxi_readdata_tmp_valid_25 <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_outstanding_wcount <= 0;
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= 0;
      _maxi_read_op_sel <= 0;
      _maxi_read_global_addr <= 0;
      _maxi_read_global_size <= 0;
      _maxi_read_local_addr <= 0;
      _maxi_read_local_stride <= 0;
      _maxi_read_local_size <= 0;
      _maxi_read_local_blocksize <= 0;
      _maxi_read_req_busy <= 0;
      _maxi_read_cur_global_size <= 0;
      _maxi_read_data_busy <= 0;
      _maxi_read_op_sel_buf <= 0;
      _maxi_read_local_addr_buf <= 0;
      _maxi_read_local_stride_buf <= 0;
      _maxi_read_local_size_buf <= 0;
      _maxi_read_local_blocksize_buf <= 0;
      _maxi_write_op_sel <= 0;
      _maxi_write_global_addr <= 0;
      _maxi_write_global_size <= 0;
      _maxi_write_local_addr <= 0;
      _maxi_write_local_stride <= 0;
      _maxi_write_local_size <= 0;
      _maxi_write_local_blocksize <= 0;
      _maxi_write_req_busy <= 0;
      _maxi_write_cur_global_size <= 0;
      _maxi_write_data_busy <= 0;
      _maxi_write_op_sel_buf <= 0;
      _maxi_write_local_addr_buf <= 0;
      _maxi_write_local_stride_buf <= 0;
      _maxi_write_size_buf <= 0;
      _maxi_write_local_blocksize_buf <= 0;
    end else begin
      if(maxi_awvalid && maxi_awready && !(maxi_bvalid && maxi_bready) && (_maxi_outstanding_wcount < 7)) begin
        _maxi_outstanding_wcount <= _maxi_outstanding_wcount + 1;
      end 
      if(!(maxi_awvalid && maxi_awready) && (maxi_bvalid && maxi_bready) && (_maxi_outstanding_wcount > 0)) begin
        _maxi_outstanding_wcount <= _maxi_outstanding_wcount - 1;
      end 
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= _saxi_register_32;
      if((control_conv2d_4 == 2) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 1;
        _maxi_read_global_addr <= mask_addr_masked_58;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_56;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_56;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_req_fsm == 0) && _maxi_read_start) begin
        _maxi_read_req_busy <= 1;
      end 
      if(_maxi_read_start && _maxi_read_req_fifo_almost_full) begin
        _maxi_read_start <= 1;
      end 
      if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && (_maxi_read_global_size <= 256) && ((mask_addr_masked_68 & 4095) + (_maxi_read_global_size << 2) >= 4096)) begin
        _maxi_read_cur_global_size <= 4096 - (mask_addr_masked_70 & 4095) >> 2;
        _maxi_read_global_size <= _maxi_read_global_size - (4096 - (mask_addr_masked_72 & 4095) >> 2);
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && (_maxi_read_global_size <= 256)) begin
        _maxi_read_cur_global_size <= _maxi_read_global_size;
        _maxi_read_global_size <= 0;
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && ((mask_addr_masked_74 & 4095) + 1024 >= 4096)) begin
        _maxi_read_cur_global_size <= 4096 - (mask_addr_masked_76 & 4095) >> 2;
        _maxi_read_global_size <= _maxi_read_global_size - (4096 - (mask_addr_masked_78 & 4095) >> 2);
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full) begin
        _maxi_read_cur_global_size <= 256;
        _maxi_read_global_size <= _maxi_read_global_size - 256;
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid)) begin
        _maxi_read_global_addr <= _maxi_read_global_addr + (_maxi_read_cur_global_size << 2);
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid) && (_maxi_read_global_size == 0)) begin
        _maxi_read_req_busy <= 0;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 4) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 2;
        _maxi_read_global_addr <= mask_addr_masked_91;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_89;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_89;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 3;
        _maxi_read_global_addr <= mask_addr_masked_107;
        _maxi_read_global_size <= _dma_write_block_local_size_102;
        _maxi_read_local_addr <= conv2d_4_filter_page_dma_offset;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_write_block_local_size_102;
        _maxi_read_local_blocksize <= _dma_read_block_local_blocksize_105;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 14) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 4;
        _maxi_read_global_addr <= mask_addr_masked_209;
        _maxi_read_global_size <= _dma_write_block_local_size_204;
        _maxi_read_local_addr <= conv2d_4_act_page_dma_offset_0;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_write_block_local_size_204;
        _maxi_read_local_blocksize <= _dma_read_block_local_blocksize_207;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 17) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 5;
        _maxi_read_global_addr <= mask_addr_masked_251;
        _maxi_read_global_size <= _dma_write_block_local_size_246;
        _maxi_read_local_addr <= conv2d_4_act_page_dma_offset_1;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_write_block_local_size_246;
        _maxi_read_local_blocksize <= _dma_read_block_local_blocksize_249;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 20) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 6;
        _maxi_read_global_addr <= mask_addr_masked_293;
        _maxi_read_global_size <= _dma_write_block_local_size_288;
        _maxi_read_local_addr <= conv2d_4_act_page_dma_offset_2;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_write_block_local_size_288;
        _maxi_read_local_blocksize <= _dma_read_block_local_blocksize_291;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 29) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 1;
        _maxi_write_global_addr <= mask_addr_masked_1137;
        _maxi_write_global_size <= _dma_write_packed_local_packed_size_1135;
        _maxi_write_local_addr <= conv2d_4_out_laddr_offset + conv2d_4_out_page_dma_offset;
        _maxi_write_local_stride <= 2;
        _maxi_write_local_size <= _dma_write_packed_local_packed_size_1135;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_req_fsm == 0) && _maxi_write_start) begin
        _maxi_write_req_busy <= 1;
      end 
      if(_maxi_write_start && _maxi_write_req_fifo_almost_full) begin
        _maxi_write_start <= 1;
      end 
      if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && (_maxi_write_global_size <= 256) && ((mask_addr_masked_1147 & 4095) + (_maxi_write_global_size << 2) >= 4096)) begin
        _maxi_write_cur_global_size <= 4096 - (mask_addr_masked_1149 & 4095) >> 2;
        _maxi_write_global_size <= _maxi_write_global_size - (4096 - (mask_addr_masked_1151 & 4095) >> 2);
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && (_maxi_write_global_size <= 256)) begin
        _maxi_write_cur_global_size <= _maxi_write_global_size;
        _maxi_write_global_size <= 0;
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && ((mask_addr_masked_1153 & 4095) + 1024 >= 4096)) begin
        _maxi_write_cur_global_size <= 4096 - (mask_addr_masked_1155 & 4095) >> 2;
        _maxi_write_global_size <= _maxi_write_global_size - (4096 - (mask_addr_masked_1157 & 4095) >> 2);
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full) begin
        _maxi_write_cur_global_size <= 256;
        _maxi_write_global_size <= _maxi_write_global_size - 256;
      end 
      if((_maxi_write_req_fsm == 1) && ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))) begin
        _maxi_write_global_addr <= _maxi_write_global_addr + (_maxi_write_cur_global_size << 2);
      end 
      if((_maxi_write_req_fsm == 1) && ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) && (_maxi_write_global_size == 0)) begin
        _maxi_write_req_busy <= 0;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_packed_rvalid_1169 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 1) && read_burst_packed_rvalid_1169 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_packed_rlast_1170) begin
        _maxi_write_data_busy <= 0;
      end 
      if((control_max_pool_serial_6 == 5) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 7;
        _maxi_read_global_addr <= mask_addr_masked_1181;
        _maxi_read_global_size <= cparam_max_pool_serial_6_act_read_size;
        _maxi_read_local_addr <= max_pool_serial_6_act_page_dma_offset;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_max_pool_serial_6_act_read_size;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_max_pool_serial_6 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 7;
        _maxi_read_global_addr <= mask_addr_masked_1187;
        _maxi_read_global_size <= cparam_max_pool_serial_6_act_read_size;
        _maxi_read_local_addr <= max_pool_serial_6_act_page_dma_offset + cparam_max_pool_serial_6_act_read_size;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_max_pool_serial_6_act_read_size;
        _maxi_read_local_blocksize <= 1;
      end 
      if((control_max_pool_serial_6 == 15) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 2;
        _maxi_write_global_addr <= mask_addr_masked_1297;
        _maxi_write_global_size <= cparam_max_pool_serial_6_out_write_size;
        _maxi_write_local_addr <= max_pool_serial_6_out_page_dma_offset;
        _maxi_write_local_stride <= 1;
        _maxi_write_local_size <= cparam_max_pool_serial_6_out_write_size;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_rvalid_1301 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 2) && read_burst_rvalid_1301 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_rlast_1302) begin
        _maxi_write_data_busy <= 0;
      end 
      if((control_matmul_23 == 2) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 8;
        _maxi_read_global_addr <= mask_addr_masked_1310;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1308;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1308;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_23 == 4) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 9;
        _maxi_read_global_addr <= mask_addr_masked_1323;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1321;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1321;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_23 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 10;
        _maxi_read_global_addr <= mask_addr_masked_1336;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1334;
        _maxi_read_local_addr <= matmul_23_filter_page_dma_offset;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1334;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 10))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_23 == 14) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 11;
        _maxi_read_global_addr <= mask_addr_masked_1349;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1347;
        _maxi_read_local_addr <= matmul_23_act_page_dma_offset_0;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1347;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 11))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_23 == 23) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 1;
        _maxi_write_global_addr <= mask_addr_masked_1633;
        _maxi_write_global_size <= _dma_write_packed_local_packed_size_1631;
        _maxi_write_local_addr <= matmul_23_out_laddr_offset + matmul_23_out_page_dma_offset;
        _maxi_write_local_stride <= 2;
        _maxi_write_local_size <= _dma_write_packed_local_packed_size_1631;
        _maxi_write_local_blocksize <= 1;
      end 
      if((control_matmul_33 == 2) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 12;
        _maxi_read_global_addr <= mask_addr_masked_1635;
        _maxi_read_global_size <= cparam_matmul_33_bias_num;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_matmul_33_bias_num;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 12))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_33 == 4) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 13;
        _maxi_read_global_addr <= mask_addr_masked_1641;
        _maxi_read_global_size <= cparam_matmul_33_scale_num;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_matmul_33_scale_num;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 13))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_33 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 14;
        _maxi_read_global_addr <= mask_addr_masked_1647;
        _maxi_read_global_size <= cparam_matmul_33_filter_read_size;
        _maxi_read_local_addr <= matmul_33_filter_page_dma_offset;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_matmul_33_filter_read_size;
        _maxi_read_local_blocksize <= cparam_matmul_33_filter_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 14))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_33 == 14) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 15;
        _maxi_read_global_addr <= mask_addr_masked_1665;
        _maxi_read_global_size <= cparam_matmul_33_act_read_size;
        _maxi_read_local_addr <= matmul_33_act_page_dma_offset_0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_matmul_33_act_read_size;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 15))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_33 == 23) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 3;
        _maxi_write_global_addr <= mask_addr_masked_2008;
        _maxi_write_global_size <= matmul_33_next_out_write_size;
        _maxi_write_local_addr <= matmul_33_out_laddr_offset + matmul_33_out_page_dma_offset;
        _maxi_write_local_stride <= 1;
        _maxi_write_local_size <= matmul_33_next_out_write_size;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_rvalid_2012 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 3) && read_burst_rvalid_2012 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_rlast_2013) begin
        _maxi_write_data_busy <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      count__maxi_read_req_fifo <= 0;
      __tmp_66_1 <= 0;
    end else begin
      if(_maxi_read_req_fifo_enq && !_maxi_read_req_fifo_full && (_maxi_read_req_fifo_deq && !_maxi_read_req_fifo_empty)) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo;
      end else if(_maxi_read_req_fifo_enq && !_maxi_read_req_fifo_full) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo + 1;
      end else if(_maxi_read_req_fifo_deq && !_maxi_read_req_fifo_empty) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo - 1;
      end 
      __tmp_66_1 <= _tmp_66;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      count__maxi_write_req_fifo <= 0;
      __tmp_1145_1 <= 0;
      __tmp_1165_1 <= 0;
    end else begin
      if(_maxi_write_req_fifo_enq && !_maxi_write_req_fifo_full && (_maxi_write_req_fifo_deq && !_maxi_write_req_fifo_empty)) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo;
      end else if(_maxi_write_req_fifo_enq && !_maxi_write_req_fifo_full) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo + 1;
      end else if(_maxi_write_req_fifo_deq && !_maxi_write_req_fifo_empty) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo - 1;
      end 
      __tmp_1145_1 <= _tmp_1145;
      __tmp_1165_1 <= _tmp_1165;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      saxi_rdata <= 0;
      saxi_rvalid <= 0;
      _saxi_rdata_cond_0_1 <= 0;
    end else begin
      if(_saxi_rdata_cond_0_1) begin
        saxi_rvalid <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid)) begin
        saxi_rdata <= axislite_rdata_46;
        saxi_rvalid <= 1;
      end 
      _saxi_rdata_cond_0_1 <= 1;
      if(saxi_rvalid && !saxi_rready) begin
        saxi_rvalid <= saxi_rvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      saxi_bvalid <= 0;
      prev_awvalid_43 <= 0;
      prev_arvalid_44 <= 0;
      writevalid_41 <= 0;
      readvalid_42 <= 0;
      addr_40 <= 0;
      _saxi_register_0 <= 0;
      _saxi_flag_0 <= 0;
      _saxi_register_1 <= 0;
      _saxi_flag_1 <= 0;
      _saxi_register_2 <= 0;
      _saxi_flag_2 <= 0;
      _saxi_register_3 <= 0;
      _saxi_flag_3 <= 0;
      _saxi_register_4 <= 0;
      _saxi_flag_4 <= 0;
      _saxi_register_5 <= 0;
      _saxi_flag_5 <= 0;
      _saxi_register_6 <= 0;
      _saxi_flag_6 <= 0;
      _saxi_register_7 <= 0;
      _saxi_flag_7 <= 0;
      _saxi_register_8 <= 0;
      _saxi_flag_8 <= 0;
      _saxi_register_9 <= 0;
      _saxi_flag_9 <= 0;
      _saxi_register_10 <= 0;
      _saxi_flag_10 <= 0;
      _saxi_register_11 <= 0;
      _saxi_flag_11 <= 0;
      _saxi_register_12 <= 0;
      _saxi_flag_12 <= 0;
      _saxi_register_13 <= 0;
      _saxi_flag_13 <= 0;
      _saxi_register_14 <= 0;
      _saxi_flag_14 <= 0;
      _saxi_register_15 <= 0;
      _saxi_flag_15 <= 0;
      _saxi_register_16 <= 0;
      _saxi_flag_16 <= 0;
      _saxi_register_17 <= 0;
      _saxi_flag_17 <= 0;
      _saxi_register_18 <= 0;
      _saxi_flag_18 <= 0;
      _saxi_register_19 <= 0;
      _saxi_flag_19 <= 0;
      _saxi_register_20 <= 0;
      _saxi_flag_20 <= 0;
      _saxi_register_21 <= 0;
      _saxi_flag_21 <= 0;
      _saxi_register_22 <= 0;
      _saxi_flag_22 <= 0;
      _saxi_register_23 <= 0;
      _saxi_flag_23 <= 0;
      _saxi_register_24 <= 0;
      _saxi_flag_24 <= 0;
      _saxi_register_25 <= 0;
      _saxi_flag_25 <= 0;
      _saxi_register_26 <= 0;
      _saxi_flag_26 <= 0;
      _saxi_register_27 <= 0;
      _saxi_flag_27 <= 0;
      _saxi_register_28 <= 0;
      _saxi_flag_28 <= 0;
      _saxi_register_29 <= 0;
      _saxi_flag_29 <= 0;
      _saxi_register_30 <= 0;
      _saxi_flag_30 <= 0;
      _saxi_register_31 <= 10495424;
      _saxi_flag_31 <= 0;
      _saxi_register_32 <= 0;
      _saxi_flag_32 <= 0;
      _saxi_register_33 <= 10205632;
      _saxi_flag_33 <= 0;
      _saxi_register_34 <= 0;
      _saxi_flag_34 <= 0;
      _saxi_register_35 <= 64;
      _saxi_flag_35 <= 0;
      _saxi_register_36 <= 8256;
      _saxi_flag_36 <= 0;
      _saxi_register_11[0] <= (0 >> 0) & 1'd1;
      _saxi_register_9[0] <= (0 >> 0) & 1'd1;
      _saxi_register_11[1] <= (0 >> 1) & 1'd1;
      _saxi_register_9[1] <= (0 >> 1) & 1'd1;
      _saxi_register_11[2] <= (0 >> 2) & 1'd1;
      _saxi_register_9[2] <= (0 >> 2) & 1'd1;
      _saxi_register_11[3] <= (0 >> 3) & 1'd1;
      _saxi_register_9[3] <= (0 >> 3) & 1'd1;
      _saxi_register_11[4] <= (0 >> 4) & 1'd1;
      _saxi_register_9[4] <= (0 >> 4) & 1'd1;
      _saxi_register_11[5] <= (0 >> 5) & 1'd1;
      _saxi_register_9[5] <= (0 >> 5) & 1'd1;
      _saxi_register_11[6] <= (0 >> 6) & 1'd1;
      _saxi_register_9[6] <= (0 >> 6) & 1'd1;
      _saxi_register_11[7] <= (0 >> 7) & 1'd1;
      _saxi_register_9[7] <= (0 >> 7) & 1'd1;
      _saxi_register_11[8] <= (0 >> 8) & 1'd1;
      _saxi_register_9[8] <= (0 >> 8) & 1'd1;
      _saxi_register_11[9] <= (0 >> 9) & 1'd1;
      _saxi_register_9[9] <= (0 >> 9) & 1'd1;
      _saxi_register_11[10] <= (0 >> 10) & 1'd1;
      _saxi_register_9[10] <= (0 >> 10) & 1'd1;
      _saxi_register_11[11] <= (0 >> 11) & 1'd1;
      _saxi_register_9[11] <= (0 >> 11) & 1'd1;
      _saxi_register_11[12] <= (0 >> 12) & 1'd1;
      _saxi_register_9[12] <= (0 >> 12) & 1'd1;
      _saxi_register_11[13] <= (0 >> 13) & 1'd1;
      _saxi_register_9[13] <= (0 >> 13) & 1'd1;
      _saxi_register_11[14] <= (0 >> 14) & 1'd1;
      _saxi_register_9[14] <= (0 >> 14) & 1'd1;
      _saxi_register_11[15] <= (0 >> 15) & 1'd1;
      _saxi_register_9[15] <= (0 >> 15) & 1'd1;
      _saxi_register_11[16] <= (0 >> 16) & 1'd1;
      _saxi_register_9[16] <= (0 >> 16) & 1'd1;
      _saxi_register_11[17] <= (0 >> 17) & 1'd1;
      _saxi_register_9[17] <= (0 >> 17) & 1'd1;
      _saxi_register_11[18] <= (0 >> 18) & 1'd1;
      _saxi_register_9[18] <= (0 >> 18) & 1'd1;
      _saxi_register_11[19] <= (0 >> 19) & 1'd1;
      _saxi_register_9[19] <= (0 >> 19) & 1'd1;
      _saxi_register_11[20] <= (0 >> 20) & 1'd1;
      _saxi_register_9[20] <= (0 >> 20) & 1'd1;
      _saxi_register_11[21] <= (0 >> 21) & 1'd1;
      _saxi_register_9[21] <= (0 >> 21) & 1'd1;
      _saxi_register_11[22] <= (0 >> 22) & 1'd1;
      _saxi_register_9[22] <= (0 >> 22) & 1'd1;
      _saxi_register_11[23] <= (0 >> 23) & 1'd1;
      _saxi_register_9[23] <= (0 >> 23) & 1'd1;
      _saxi_register_11[24] <= (0 >> 24) & 1'd1;
      _saxi_register_9[24] <= (0 >> 24) & 1'd1;
      _saxi_register_11[25] <= (0 >> 25) & 1'd1;
      _saxi_register_9[25] <= (0 >> 25) & 1'd1;
      _saxi_register_11[26] <= (0 >> 26) & 1'd1;
      _saxi_register_9[26] <= (0 >> 26) & 1'd1;
      _saxi_register_11[27] <= (0 >> 27) & 1'd1;
      _saxi_register_9[27] <= (0 >> 27) & 1'd1;
      _saxi_register_11[28] <= (0 >> 28) & 1'd1;
      _saxi_register_9[28] <= (0 >> 28) & 1'd1;
      _saxi_register_11[29] <= (0 >> 29) & 1'd1;
      _saxi_register_9[29] <= (0 >> 29) & 1'd1;
      _saxi_register_11[30] <= (0 >> 30) & 1'd1;
      _saxi_register_9[30] <= (0 >> 30) & 1'd1;
      _saxi_register_11[31] <= (0 >> 31) & 1'd1;
      _saxi_register_9[31] <= (0 >> 31) & 1'd1;
      internal_state_counter <= 0;
    end else begin
      if(saxi_bvalid && saxi_bready) begin
        saxi_bvalid <= 0;
      end 
      if(saxi_wvalid && saxi_wready) begin
        saxi_bvalid <= 1;
      end 
      prev_awvalid_43 <= saxi_awvalid;
      prev_arvalid_44 <= saxi_arvalid;
      writevalid_41 <= 0;
      readvalid_42 <= 0;
      if(saxi_awready && saxi_awvalid && !saxi_bvalid) begin
        addr_40 <= saxi_awaddr;
        writevalid_41 <= 1;
      end else if(saxi_arready && saxi_arvalid) begin
        addr_40 <= saxi_araddr;
        readvalid_42 <= 1;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 0)) begin
        _saxi_register_0 <= axislite_resetval_48;
        _saxi_flag_0 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 1)) begin
        _saxi_register_1 <= axislite_resetval_48;
        _saxi_flag_1 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 2)) begin
        _saxi_register_2 <= axislite_resetval_48;
        _saxi_flag_2 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 3)) begin
        _saxi_register_3 <= axislite_resetval_48;
        _saxi_flag_3 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 4)) begin
        _saxi_register_4 <= axislite_resetval_48;
        _saxi_flag_4 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 5)) begin
        _saxi_register_5 <= axislite_resetval_48;
        _saxi_flag_5 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 6)) begin
        _saxi_register_6 <= axislite_resetval_48;
        _saxi_flag_6 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 7)) begin
        _saxi_register_7 <= axislite_resetval_48;
        _saxi_flag_7 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 8)) begin
        _saxi_register_8 <= axislite_resetval_48;
        _saxi_flag_8 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 9)) begin
        _saxi_register_9 <= axislite_resetval_48;
        _saxi_flag_9 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 10)) begin
        _saxi_register_10 <= axislite_resetval_48;
        _saxi_flag_10 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 11)) begin
        _saxi_register_11 <= axislite_resetval_48;
        _saxi_flag_11 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 12)) begin
        _saxi_register_12 <= axislite_resetval_48;
        _saxi_flag_12 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 13)) begin
        _saxi_register_13 <= axislite_resetval_48;
        _saxi_flag_13 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 14)) begin
        _saxi_register_14 <= axislite_resetval_48;
        _saxi_flag_14 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 15)) begin
        _saxi_register_15 <= axislite_resetval_48;
        _saxi_flag_15 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 16)) begin
        _saxi_register_16 <= axislite_resetval_48;
        _saxi_flag_16 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 17)) begin
        _saxi_register_17 <= axislite_resetval_48;
        _saxi_flag_17 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 18)) begin
        _saxi_register_18 <= axislite_resetval_48;
        _saxi_flag_18 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 19)) begin
        _saxi_register_19 <= axislite_resetval_48;
        _saxi_flag_19 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 20)) begin
        _saxi_register_20 <= axislite_resetval_48;
        _saxi_flag_20 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 21)) begin
        _saxi_register_21 <= axislite_resetval_48;
        _saxi_flag_21 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 22)) begin
        _saxi_register_22 <= axislite_resetval_48;
        _saxi_flag_22 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 23)) begin
        _saxi_register_23 <= axislite_resetval_48;
        _saxi_flag_23 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 24)) begin
        _saxi_register_24 <= axislite_resetval_48;
        _saxi_flag_24 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 25)) begin
        _saxi_register_25 <= axislite_resetval_48;
        _saxi_flag_25 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 26)) begin
        _saxi_register_26 <= axislite_resetval_48;
        _saxi_flag_26 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 27)) begin
        _saxi_register_27 <= axislite_resetval_48;
        _saxi_flag_27 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 28)) begin
        _saxi_register_28 <= axislite_resetval_48;
        _saxi_flag_28 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 29)) begin
        _saxi_register_29 <= axislite_resetval_48;
        _saxi_flag_29 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 30)) begin
        _saxi_register_30 <= axislite_resetval_48;
        _saxi_flag_30 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 31)) begin
        _saxi_register_31 <= axislite_resetval_48;
        _saxi_flag_31 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 32)) begin
        _saxi_register_32 <= axislite_resetval_48;
        _saxi_flag_32 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 33)) begin
        _saxi_register_33 <= axislite_resetval_48;
        _saxi_flag_33 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 34)) begin
        _saxi_register_34 <= axislite_resetval_48;
        _saxi_flag_34 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 35)) begin
        _saxi_register_35 <= axislite_resetval_48;
        _saxi_flag_35 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 36)) begin
        _saxi_register_36 <= axislite_resetval_48;
        _saxi_flag_36 <= 0;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 0)) begin
        _saxi_register_0 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 1)) begin
        _saxi_register_1 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 2)) begin
        _saxi_register_2 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 3)) begin
        _saxi_register_3 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 4)) begin
        _saxi_register_4 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 5)) begin
        _saxi_register_5 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 6)) begin
        _saxi_register_6 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 7)) begin
        _saxi_register_7 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 8)) begin
        _saxi_register_8 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 9)) begin
        _saxi_register_9 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 10)) begin
        _saxi_register_10 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 11)) begin
        _saxi_register_11 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 12)) begin
        _saxi_register_12 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 13)) begin
        _saxi_register_13 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 14)) begin
        _saxi_register_14 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 15)) begin
        _saxi_register_15 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 16)) begin
        _saxi_register_16 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 17)) begin
        _saxi_register_17 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 18)) begin
        _saxi_register_18 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 19)) begin
        _saxi_register_19 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 20)) begin
        _saxi_register_20 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 21)) begin
        _saxi_register_21 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 22)) begin
        _saxi_register_22 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 23)) begin
        _saxi_register_23 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 24)) begin
        _saxi_register_24 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 25)) begin
        _saxi_register_25 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 26)) begin
        _saxi_register_26 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 27)) begin
        _saxi_register_27 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 28)) begin
        _saxi_register_28 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 29)) begin
        _saxi_register_29 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 30)) begin
        _saxi_register_30 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 31)) begin
        _saxi_register_31 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 32)) begin
        _saxi_register_32 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 33)) begin
        _saxi_register_33 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 34)) begin
        _saxi_register_34 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 35)) begin
        _saxi_register_35 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 36)) begin
        _saxi_register_36 <= saxi_wdata;
      end 
      if(_saxi_register_11[0] == 1) begin
        _saxi_register_11[0] <= 0;
        _saxi_register_9[0] <= 0;
      end 
      if(_saxi_register_11[1] == 1) begin
        _saxi_register_11[1] <= 0;
        _saxi_register_9[1] <= 0;
      end 
      if(_saxi_register_11[2] == 1) begin
        _saxi_register_11[2] <= 0;
        _saxi_register_9[2] <= 0;
      end 
      if(_saxi_register_11[3] == 1) begin
        _saxi_register_11[3] <= 0;
        _saxi_register_9[3] <= 0;
      end 
      if(_saxi_register_11[4] == 1) begin
        _saxi_register_11[4] <= 0;
        _saxi_register_9[4] <= 0;
      end 
      if(_saxi_register_11[5] == 1) begin
        _saxi_register_11[5] <= 0;
        _saxi_register_9[5] <= 0;
      end 
      if(_saxi_register_11[6] == 1) begin
        _saxi_register_11[6] <= 0;
        _saxi_register_9[6] <= 0;
      end 
      if(_saxi_register_11[7] == 1) begin
        _saxi_register_11[7] <= 0;
        _saxi_register_9[7] <= 0;
      end 
      if(_saxi_register_11[8] == 1) begin
        _saxi_register_11[8] <= 0;
        _saxi_register_9[8] <= 0;
      end 
      if(_saxi_register_11[9] == 1) begin
        _saxi_register_11[9] <= 0;
        _saxi_register_9[9] <= 0;
      end 
      if(_saxi_register_11[10] == 1) begin
        _saxi_register_11[10] <= 0;
        _saxi_register_9[10] <= 0;
      end 
      if(_saxi_register_11[11] == 1) begin
        _saxi_register_11[11] <= 0;
        _saxi_register_9[11] <= 0;
      end 
      if(_saxi_register_11[12] == 1) begin
        _saxi_register_11[12] <= 0;
        _saxi_register_9[12] <= 0;
      end 
      if(_saxi_register_11[13] == 1) begin
        _saxi_register_11[13] <= 0;
        _saxi_register_9[13] <= 0;
      end 
      if(_saxi_register_11[14] == 1) begin
        _saxi_register_11[14] <= 0;
        _saxi_register_9[14] <= 0;
      end 
      if(_saxi_register_11[15] == 1) begin
        _saxi_register_11[15] <= 0;
        _saxi_register_9[15] <= 0;
      end 
      if(_saxi_register_11[16] == 1) begin
        _saxi_register_11[16] <= 0;
        _saxi_register_9[16] <= 0;
      end 
      if(_saxi_register_11[17] == 1) begin
        _saxi_register_11[17] <= 0;
        _saxi_register_9[17] <= 0;
      end 
      if(_saxi_register_11[18] == 1) begin
        _saxi_register_11[18] <= 0;
        _saxi_register_9[18] <= 0;
      end 
      if(_saxi_register_11[19] == 1) begin
        _saxi_register_11[19] <= 0;
        _saxi_register_9[19] <= 0;
      end 
      if(_saxi_register_11[20] == 1) begin
        _saxi_register_11[20] <= 0;
        _saxi_register_9[20] <= 0;
      end 
      if(_saxi_register_11[21] == 1) begin
        _saxi_register_11[21] <= 0;
        _saxi_register_9[21] <= 0;
      end 
      if(_saxi_register_11[22] == 1) begin
        _saxi_register_11[22] <= 0;
        _saxi_register_9[22] <= 0;
      end 
      if(_saxi_register_11[23] == 1) begin
        _saxi_register_11[23] <= 0;
        _saxi_register_9[23] <= 0;
      end 
      if(_saxi_register_11[24] == 1) begin
        _saxi_register_11[24] <= 0;
        _saxi_register_9[24] <= 0;
      end 
      if(_saxi_register_11[25] == 1) begin
        _saxi_register_11[25] <= 0;
        _saxi_register_9[25] <= 0;
      end 
      if(_saxi_register_11[26] == 1) begin
        _saxi_register_11[26] <= 0;
        _saxi_register_9[26] <= 0;
      end 
      if(_saxi_register_11[27] == 1) begin
        _saxi_register_11[27] <= 0;
        _saxi_register_9[27] <= 0;
      end 
      if(_saxi_register_11[28] == 1) begin
        _saxi_register_11[28] <= 0;
        _saxi_register_9[28] <= 0;
      end 
      if(_saxi_register_11[29] == 1) begin
        _saxi_register_11[29] <= 0;
        _saxi_register_9[29] <= 0;
      end 
      if(_saxi_register_11[30] == 1) begin
        _saxi_register_11[30] <= 0;
        _saxi_register_9[30] <= 0;
      end 
      if(_saxi_register_11[31] == 1) begin
        _saxi_register_11[31] <= 0;
        _saxi_register_9[31] <= 0;
      end 
      if(irq_busy_edge_51) begin
        _saxi_register_9[0] <= irq_busy_edge_51;
      end 
      if(irq_extern_edge_53) begin
        _saxi_register_9[1] <= irq_extern_edge_53;
      end 
      if(main_fsm == 0) begin
        _saxi_register_5 <= 0;
        _saxi_register_6 <= 0;
        _saxi_register_7 <= 0;
      end 
      if(main_fsm == 1) begin
        internal_state_counter <= 0;
        _saxi_register_12 <= 0;
      end else if(main_fsm == _saxi_register_13) begin
        if(internal_state_counter == _saxi_register_14) begin
          internal_state_counter <= 0;
          _saxi_register_12 <= _saxi_register_12 + 1;
        end else begin
          internal_state_counter <= internal_state_counter + 1;
        end
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_0 <= 1;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_1 <= 1;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_2 <= 1;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_3 <= 1;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_4 <= 1;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 1) && 1) begin
        _saxi_register_5 <= 1;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_6 <= 1;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_7 <= 1;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_8 <= 1;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_9 <= 1;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_10 <= 1;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_11 <= 1;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_12 <= 1;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_13 <= 1;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_14 <= 1;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_15 <= 1;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_16 <= 1;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_17 <= 1;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_18 <= 1;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_19 <= 1;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_20 <= 1;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_21 <= 1;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_22 <= 1;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_23 <= 1;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_24 <= 1;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_25 <= 1;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_26 <= 1;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_27 <= 1;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_28 <= 1;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_29 <= 1;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_30 <= 1;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_31 <= 1;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_32 <= 1;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_33 <= 1;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_34 <= 1;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_35 <= 1;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_36 <= 1;
        _saxi_flag_36 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 2) && 1) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_14 <= 0;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_15 <= 0;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_16 <= 0;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_17 <= 0;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_18 <= 0;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_19 <= 0;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_20 <= 0;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_21 <= 0;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_22 <= 0;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_23 <= 0;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_24 <= 0;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_25 <= 0;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_26 <= 0;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_27 <= 0;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_28 <= 0;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_29 <= 0;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_30 <= 0;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_31 <= 0;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_32 <= 0;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_33 <= 0;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_34 <= 0;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_35 <= 0;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_36 <= 0;
        _saxi_flag_36 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 88) && 1) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_14 <= 0;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_15 <= 0;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_16 <= 0;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_17 <= 0;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_18 <= 0;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_19 <= 0;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_20 <= 0;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_21 <= 0;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_22 <= 0;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_23 <= 0;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_24 <= 0;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_25 <= 0;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_26 <= 0;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_27 <= 0;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_28 <= 0;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_29 <= 0;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_30 <= 0;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_31 <= 0;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_32 <= 0;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_33 <= 0;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_34 <= 0;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_35 <= 0;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 88) && 0) begin
        _saxi_register_36 <= 0;
        _saxi_flag_36 <= 0;
      end 
    end
  end

  localparam _saxi_register_fsm_1 = 1;
  localparam _saxi_register_fsm_2 = 2;
  localparam _saxi_register_fsm_3 = 3;
  localparam _saxi_register_fsm_4 = 4;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _saxi_register_fsm <= _saxi_register_fsm_init;
      axis_maskaddr_45 <= 0;
    end else begin
      case(_saxi_register_fsm)
        _saxi_register_fsm_init: begin
          if(readvalid_42 || writevalid_41) begin
            axis_maskaddr_45 <= (addr_40 >> _saxi_shift) & _saxi_mask;
          end 
          if(readvalid_42) begin
            _saxi_register_fsm <= _saxi_register_fsm_1;
          end 
          if(writevalid_41) begin
            _saxi_register_fsm <= _saxi_register_fsm_3;
          end 
        end
        _saxi_register_fsm_1: begin
          if(saxi_rready || !saxi_rvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_2;
          end 
        end
        _saxi_register_fsm_2: begin
          if(saxi_rready && saxi_rvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_init;
          end 
        end
        _saxi_register_fsm_3: begin
          if(saxi_wvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_4;
          end 
        end
        _saxi_register_fsm_4: begin
          if(saxi_bready && saxi_bvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    _rst_logic_1 <= rst_logic;
    _rst_logic_2 <= _rst_logic_1;
    RST <= rst_logic | _rst_logic_1 | _rst_logic_2;
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq <= 0;
    end else begin
      irq <= |irq_49;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq_busy_edge_50 <= 0;
    end else begin
      irq_busy_edge_50 <= irq_busy;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq_extern_edge_52 <= 0;
    end else begin
      irq_extern_edge_52 <= irq_extern;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1406_1 <= 0;
    end else begin
      __tmp_1406_1 <= _tmp_1406;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1408_1 <= 0;
    end else begin
      __tmp_1408_1 <= _tmp_1408;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1192_1 <= 0;
    end else begin
      __tmp_1192_1 <= _tmp_1192;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1397_1 <= 0;
    end else begin
      __tmp_1397_1 <= _tmp_1397;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1399_1 <= 0;
    end else begin
      __tmp_1399_1 <= _tmp_1399;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1304_1 <= 0;
      __tmp_1701_1 <= 0;
    end else begin
      __tmp_1304_1 <= _tmp_1304;
      __tmp_1701_1 <= _tmp_1701;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1695_1 <= 0;
    end else begin
      __tmp_1695_1 <= _tmp_1695;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1698_1 <= 0;
    end else begin
      __tmp_1698_1 <= _tmp_1698;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_367_1 <= 0;
      __tmp_1368_1 <= 0;
    end else begin
      __tmp_367_1 <= _tmp_367;
      __tmp_1368_1 <= _tmp_1368;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_369_1 <= 0;
      __tmp_1370_1 <= 0;
    end else begin
      __tmp_369_1 <= _tmp_369;
      __tmp_1370_1 <= _tmp_1370;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_376_1 <= 0;
      __tmp_1378_1 <= 0;
    end else begin
      __tmp_376_1 <= _tmp_376;
      __tmp_1378_1 <= _tmp_1378;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_378_1 <= 0;
      __tmp_1380_1 <= 0;
    end else begin
      __tmp_378_1 <= _tmp_378;
      __tmp_1380_1 <= _tmp_1380;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_385_1 <= 0;
    end else begin
      __tmp_385_1 <= _tmp_385;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_387_1 <= 0;
    end else begin
      __tmp_387_1 <= _tmp_387;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_394_1 <= 0;
    end else begin
      __tmp_394_1 <= _tmp_394;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_396_1 <= 0;
    end else begin
      __tmp_396_1 <= _tmp_396;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_403_1 <= 0;
    end else begin
      __tmp_403_1 <= _tmp_403;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_405_1 <= 0;
    end else begin
      __tmp_405_1 <= _tmp_405;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_412_1 <= 0;
    end else begin
      __tmp_412_1 <= _tmp_412;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_414_1 <= 0;
    end else begin
      __tmp_414_1 <= _tmp_414;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_421_1 <= 0;
    end else begin
      __tmp_421_1 <= _tmp_421;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_423_1 <= 0;
    end else begin
      __tmp_423_1 <= _tmp_423;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_430_1 <= 0;
    end else begin
      __tmp_430_1 <= _tmp_430;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_432_1 <= 0;
    end else begin
      __tmp_432_1 <= _tmp_432;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_439_1 <= 0;
    end else begin
      __tmp_439_1 <= _tmp_439;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_441_1 <= 0;
    end else begin
      __tmp_441_1 <= _tmp_441;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1173_1 <= 0;
    end else begin
      __tmp_1173_1 <= _tmp_1173;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1177_1 <= 0;
    end else begin
      __tmp_1177_1 <= _tmp_1177;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_338_1 <= 0;
    end else begin
      __tmp_338_1 <= _tmp_338;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_340_1 <= 0;
    end else begin
      __tmp_340_1 <= _tmp_340;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_348_1 <= 0;
    end else begin
      __tmp_348_1 <= _tmp_348;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_350_1 <= 0;
    end else begin
      __tmp_350_1 <= _tmp_350;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_448_1 <= 0;
    end else begin
      __tmp_448_1 <= _tmp_448;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_450_1 <= 0;
    end else begin
      __tmp_450_1 <= _tmp_450;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_457_1 <= 0;
    end else begin
      __tmp_457_1 <= _tmp_457;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_459_1 <= 0;
    end else begin
      __tmp_459_1 <= _tmp_459;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_466_1 <= 0;
    end else begin
      __tmp_466_1 <= _tmp_466;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_468_1 <= 0;
    end else begin
      __tmp_468_1 <= _tmp_468;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_475_1 <= 0;
    end else begin
      __tmp_475_1 <= _tmp_475;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_477_1 <= 0;
    end else begin
      __tmp_477_1 <= _tmp_477;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_484_1 <= 0;
    end else begin
      __tmp_484_1 <= _tmp_484;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_486_1 <= 0;
    end else begin
      __tmp_486_1 <= _tmp_486;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_493_1 <= 0;
    end else begin
      __tmp_493_1 <= _tmp_493;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_495_1 <= 0;
    end else begin
      __tmp_495_1 <= _tmp_495;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_502_1 <= 0;
    end else begin
      __tmp_502_1 <= _tmp_502;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_504_1 <= 0;
    end else begin
      __tmp_504_1 <= _tmp_504;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_511_1 <= 0;
    end else begin
      __tmp_511_1 <= _tmp_511;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_513_1 <= 0;
    end else begin
      __tmp_513_1 <= _tmp_513;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_520_1 <= 0;
    end else begin
      __tmp_520_1 <= _tmp_520;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_522_1 <= 0;
    end else begin
      __tmp_522_1 <= _tmp_522;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_2015_1 <= 0;
    end else begin
      __tmp_2015_1 <= _tmp_2015;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1678_1 <= 0;
    end else begin
      __tmp_1678_1 <= _tmp_1678;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1682_1 <= 0;
    end else begin
      __tmp_1682_1 <= _tmp_1682;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _acc_0_x_source_ram_renable <= 0;
      _acc_0_x_source_fifo_deq <= 0;
      _acc_0_x_idle <= 1;
      _acc_0_rshift_source_ram_renable <= 0;
      _acc_0_rshift_source_fifo_deq <= 0;
      _acc_0_rshift_idle <= 1;
      _acc_0_sum_sink_wenable <= 0;
      _acc_0_sum_sink_fifo_enq <= 0;
      _acc_0_valid_sink_wenable <= 0;
      _acc_0_valid_sink_fifo_enq <= 0;
      __acc_0_stream_ivalid_1 <= 0;
      __acc_0_stream_ivalid_2 <= 0;
      __acc_0_stream_ivalid_3 <= 0;
      __acc_0_stream_ivalid_4 <= 0;
      __acc_0_stream_ivalid_5 <= 0;
      _greaterthan_data_3 <= 0;
      _minus_data_5 <= 0;
      _reduceadd_data_16 <= 1'sd0;
      _reduceadd_count_16 <= 0;
      _reduceadd_prev_count_max_16 <= 0;
      _pulse_data_18 <= 1'sd0;
      _pulse_count_18 <= 0;
      _pulse_prev_count_max_18 <= 0;
      __delay_data_894__variable_1 <= 0;
      _sll_data_7 <= 0;
      __delay_data_891_greaterthan_3 <= 0;
      __delay_data_892_reduceadd_16 <= 0;
      __delay_data_895__delay_894__variable_1 <= 0;
      __delay_data_898_pulse_18 <= 0;
      _cond_data_13 <= 0;
      __delay_data_893__delay_892_reduceadd_16 <= 0;
      __delay_data_896__delay_895__delay_894__variable_1 <= 0;
      __delay_data_899__delay_898_pulse_18 <= 0;
      _plus_data_20 <= 0;
      __delay_data_897__delay_896__delay_895__delay_894__variable_1 <= 0;
      __delay_data_900__delay_899__delay_898_pulse_18 <= 0;
      _sra_data_21 <= 0;
      __delay_data_901__delay_900__delay_899__delay_898_pulse_18 <= 0;
      __variable_wdata_15 <= 0;
      __variable_wdata_0 <= 0;
      __variable_wdata_1 <= 0;
      __variable_wdata_2 <= 0;
      _tmp_951 <= 0;
      _tmp_952 <= 0;
      _tmp_953 <= 0;
      _tmp_954 <= 0;
      _tmp_955 <= 0;
      _tmp_956 <= 0;
      _tmp_957 <= 0;
      _tmp_958 <= 0;
      _tmp_959 <= 0;
      _tmp_960 <= 0;
      _tmp_961 <= 0;
      _tmp_962 <= 0;
      _tmp_963 <= 0;
      _tmp_964 <= 0;
      _tmp_965 <= 0;
      _tmp_966 <= 0;
      _tmp_967 <= 0;
      _tmp_968 <= 0;
      _tmp_969 <= 0;
      _tmp_970 <= 0;
      _tmp_971 <= 0;
      _tmp_972 <= 0;
      _tmp_973 <= 0;
      _tmp_974 <= 0;
      _tmp_975 <= 0;
      _tmp_976 <= 0;
      _tmp_977 <= 0;
      _tmp_978 <= 0;
      _tmp_979 <= 0;
      _tmp_980 <= 0;
      _tmp_981 <= 0;
      _tmp_982 <= 0;
      _acc_0_busy_reg <= 0;
    end else begin
      if(_acc_0_stream_oready) begin
        _acc_0_x_source_ram_renable <= 0;
        _acc_0_x_source_fifo_deq <= 0;
      end 
      _acc_0_x_idle <= _acc_0_x_idle;
      if(_acc_0_stream_oready) begin
        _acc_0_rshift_source_ram_renable <= 0;
        _acc_0_rshift_source_fifo_deq <= 0;
      end 
      _acc_0_rshift_idle <= _acc_0_rshift_idle;
      if(_acc_0_stream_oready) begin
        _acc_0_sum_sink_wenable <= 0;
        _acc_0_sum_sink_fifo_enq <= 0;
      end 
      if(_acc_0_stream_oready) begin
        _acc_0_valid_sink_wenable <= 0;
        _acc_0_valid_sink_fifo_enq <= 0;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_1 <= _acc_0_stream_ivalid;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_2 <= __acc_0_stream_ivalid_1;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_3 <= __acc_0_stream_ivalid_2;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_4 <= __acc_0_stream_ivalid_3;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_5 <= __acc_0_stream_ivalid_4;
      end 
      if(_acc_0_stream_oready) begin
        _greaterthan_data_3 <= acc_0_rshift_data > 1'sd0;
      end 
      if(_acc_0_stream_oready) begin
        _minus_data_5 <= acc_0_rshift_data - 2'sd1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready && _reduceadd_reset_cond_16) begin
        _reduceadd_data_16 <= 1'sd0;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _reduceadd_count_16 <= (_reduceadd_current_count_16 >= acc_0_size_data - 1)? 0 : _reduceadd_current_count_16 + 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _reduceadd_prev_count_max_16 <= _reduceadd_current_count_16 >= acc_0_size_data - 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _reduceadd_data_16 <= _reduceadd_current_data_16 + acc_0_x_data;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready && _pulse_reset_cond_18) begin
        _pulse_data_18 <= 1'sd0;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _pulse_count_18 <= (_pulse_current_count_18 >= acc_0_size_data - 1)? 0 : _pulse_current_count_18 + 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _pulse_prev_count_max_18 <= _pulse_current_count_18 >= acc_0_size_data - 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _pulse_data_18 <= _pulse_current_count_18 >= acc_0_size_data - 1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_894__variable_1 <= acc_0_rshift_data;
      end 
      if(_acc_0_stream_oready) begin
        _sll_data_7 <= 2'sd1 << _minus_data_5;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_891_greaterthan_3 <= _greaterthan_data_3;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_892_reduceadd_16 <= _reduceadd_data_16;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_895__delay_894__variable_1 <= __delay_data_894__variable_1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_898_pulse_18 <= _pulse_data_18;
      end 
      if(_acc_0_stream_oready) begin
        _cond_data_13 <= (__delay_data_891_greaterthan_3)? _sll_data_7 : 1'sd0;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_893__delay_892_reduceadd_16 <= __delay_data_892_reduceadd_16;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_896__delay_895__delay_894__variable_1 <= __delay_data_895__delay_894__variable_1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_899__delay_898_pulse_18 <= __delay_data_898_pulse_18;
      end 
      if(_acc_0_stream_oready) begin
        _plus_data_20 <= __delay_data_893__delay_892_reduceadd_16 + _cond_data_13;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_897__delay_896__delay_895__delay_894__variable_1 <= __delay_data_896__delay_895__delay_894__variable_1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_900__delay_899__delay_898_pulse_18 <= __delay_data_899__delay_898_pulse_18;
      end 
      if(_acc_0_stream_oready) begin
        _sra_data_21 <= _plus_data_20 >>> __delay_data_897__delay_896__delay_895__delay_894__variable_1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_901__delay_900__delay_899__delay_898_pulse_18 <= __delay_data_900__delay_899__delay_898_pulse_18;
      end 
      if(__stream_conv2d_4_stream_ivalid_13 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_15 <= __delay_data_1293__delay_1292__delay_1291____variable_344;
      end 
      if(__stream_conv2d_4_stream_ivalid_13 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_0 <= __substreamoutput_data_889;
      end 
      if(__stream_conv2d_4_stream_ivalid_13 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1 <= __delay_data_1305__delay_1304__delay_1303__delay_1302___plus_902;
      end 
      if(__stream_conv2d_4_stream_ivalid_13 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_2 <= __delay_data_1318__delay_1317__delay_1316____variable_339;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_951 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_952 <= _tmp_951;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_953 <= _tmp_952;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_954 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_955 <= _tmp_954;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_956 <= _tmp_955;
      end 
      if(_acc_0_stream_oready && _tmp_956) begin
        __variable_wdata_15 <= 1;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_957 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_958 <= _tmp_957;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_959 <= _tmp_958;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_960 <= _tmp_959;
      end 
      if(_acc_0_stream_oready && _tmp_960) begin
        __variable_wdata_15 <= 0;
      end 
      if(_acc_0_stream_oready && 1'd0) begin
        __variable_wdata_15 <= 1;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_961 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_962 <= _tmp_961;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_963 <= _tmp_962;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_964 <= _tmp_963;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_965 <= _tmp_964;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_966 <= _tmp_965;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_967 <= _tmp_966;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_968 <= _acc_0_source_stop;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_969 <= _tmp_968;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_970 <= _tmp_969;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_971 <= _tmp_970;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_972 <= _tmp_971;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_973 <= _tmp_972;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_974 <= _tmp_973;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_975 <= _acc_0_source_busy;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_976 <= _tmp_975;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_977 <= _tmp_976;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_978 <= _tmp_977;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_979 <= _tmp_978;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_980 <= _tmp_979;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_981 <= _tmp_980;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_982 <= _acc_0_sink_busy;
      end 
      if(!_acc_0_sink_busy && _tmp_982) begin
        _acc_0_busy_reg <= 0;
      end 
      if(_acc_0_source_busy) begin
        _acc_0_busy_reg <= 1;
      end 
      if(__stream_matmul_23_stream_ivalid_11 && _stream_matmul_23_stream_oready) begin
        __variable_wdata_15 <= __delay_data_1414__delay_1413__delay_1412____variable_961;
      end 
      if(__stream_matmul_23_stream_ivalid_11 && _stream_matmul_23_stream_oready) begin
        __variable_wdata_0 <= __substreamoutput_data_1038;
      end 
      if(__stream_matmul_23_stream_ivalid_11 && _stream_matmul_23_stream_oready) begin
        __variable_wdata_1 <= __delay_data_1424__delay_1423__delay_1422___plus_1040;
      end 
      if(__stream_matmul_23_stream_ivalid_11 && _stream_matmul_23_stream_oready) begin
        __variable_wdata_2 <= __delay_data_1435__delay_1434__delay_1433____variable_956;
      end 
      if(__stream_matmul_33_stream_ivalid_14 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_15 <= __delay_data_1536__delay_1535__delay_1534____variable_1057;
      end 
      if(__stream_matmul_33_stream_ivalid_14 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_0 <= __substreamoutput_data_1197;
      end 
      if(__stream_matmul_33_stream_ivalid_14 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_1 <= __delay_data_1549__delay_1548__delay_1547___plus_1199;
      end 
      if(__stream_matmul_33_stream_ivalid_14 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_2 <= __delay_data_1563__delay_1562__delay_1561____variable_1052;
      end 
    end
  end

  localparam _acc_0_fsm_1 = 1;
  localparam _acc_0_fsm_2 = 2;
  localparam _acc_0_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _acc_0_fsm <= _acc_0_fsm_init;
      _acc_0_source_start <= 0;
      _acc_0_source_busy <= 0;
      _acc_0_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_13 && _stream_conv2d_4_stream_oready) begin
        _acc_0_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _acc_0_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_acc_0_stream_oready && _tmp_953) begin
        _acc_0_stream_ivalid <= 1;
      end 
      if(_acc_0_stream_oready && 1'd0) begin
        _acc_0_stream_ivalid <= 0;
      end 
      if(__stream_matmul_23_stream_ivalid_11 && _stream_matmul_23_stream_oready) begin
        _acc_0_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_23_stream_oready && _stream_matmul_23_busy) begin
        _acc_0_source_busy <= _stream_matmul_23_source_busy;
      end 
      if(__stream_matmul_33_stream_ivalid_14 && _stream_matmul_33_stream_oready) begin
        _acc_0_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_busy) begin
        _acc_0_source_busy <= _stream_matmul_33_source_busy;
      end 
      case(_acc_0_fsm)
        _acc_0_fsm_init: begin
          if(_acc_0_run_flag) begin
            _acc_0_source_start <= 1;
          end 
          if(_acc_0_run_flag) begin
            _acc_0_fsm <= _acc_0_fsm_1;
          end 
        end
        _acc_0_fsm_1: begin
          if(_acc_0_source_start && _acc_0_stream_oready) begin
            _acc_0_source_start <= 0;
            _acc_0_source_busy <= 1;
          end 
          if(_acc_0_source_start && _acc_0_stream_oready) begin
            _acc_0_fsm <= _acc_0_fsm_2;
          end 
        end
        _acc_0_fsm_2: begin
          if(_acc_0_stream_oready) begin
            _acc_0_fsm <= _acc_0_fsm_3;
          end 
        end
        _acc_0_fsm_3: begin
          if(_acc_0_stream_oready && 1'd0) begin
            _acc_0_source_busy <= 0;
          end 
          if(_acc_0_stream_oready && 1'd0 && _acc_0_run_flag) begin
            _acc_0_source_start <= 1;
          end 
          if(_acc_0_stream_oready && 1'd0) begin
            _acc_0_fsm <= _acc_0_fsm_init;
          end 
          if(_acc_0_stream_oready && 1'd0 && _acc_0_run_flag) begin
            _acc_0_fsm <= _acc_0_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _acc_1_x_source_ram_renable <= 0;
      _acc_1_x_source_fifo_deq <= 0;
      _acc_1_x_idle <= 1;
      _acc_1_rshift_source_ram_renable <= 0;
      _acc_1_rshift_source_fifo_deq <= 0;
      _acc_1_rshift_idle <= 1;
      _acc_1_sum_sink_wenable <= 0;
      _acc_1_sum_sink_fifo_enq <= 0;
      _acc_1_valid_sink_wenable <= 0;
      _acc_1_valid_sink_fifo_enq <= 0;
      __acc_1_stream_ivalid_1 <= 0;
      __acc_1_stream_ivalid_2 <= 0;
      __acc_1_stream_ivalid_3 <= 0;
      __acc_1_stream_ivalid_4 <= 0;
      __acc_1_stream_ivalid_5 <= 0;
      _greaterthan_data_25 <= 0;
      _minus_data_27 <= 0;
      _reduceadd_data_38 <= 1'sd0;
      _reduceadd_count_38 <= 0;
      _reduceadd_prev_count_max_38 <= 0;
      _pulse_data_40 <= 1'sd0;
      _pulse_count_40 <= 0;
      _pulse_prev_count_max_40 <= 0;
      __delay_data_1223__variable_23 <= 0;
      _sll_data_29 <= 0;
      __delay_data_1220_greaterthan_25 <= 0;
      __delay_data_1221_reduceadd_38 <= 0;
      __delay_data_1224__delay_1223__variable_23 <= 0;
      __delay_data_1227_pulse_40 <= 0;
      _cond_data_35 <= 0;
      __delay_data_1222__delay_1221_reduceadd_38 <= 0;
      __delay_data_1225__delay_1224__delay_1223__variable_23 <= 0;
      __delay_data_1228__delay_1227_pulse_40 <= 0;
      _plus_data_42 <= 0;
      __delay_data_1226__delay_1225__delay_1224____variable_23 <= 0;
      __delay_data_1229__delay_1228__delay_1227_pulse_40 <= 0;
      _sra_data_43 <= 0;
      __delay_data_1230__delay_1229__delay_1228__delay_1227_pulse_40 <= 0;
      __variable_wdata_37 <= 0;
      __variable_wdata_22 <= 0;
      __variable_wdata_23 <= 0;
      __variable_wdata_24 <= 0;
      _tmp_1828 <= 0;
      _tmp_1829 <= 0;
      _tmp_1830 <= 0;
      _tmp_1831 <= 0;
      _tmp_1832 <= 0;
      _tmp_1833 <= 0;
      _tmp_1834 <= 0;
      _tmp_1835 <= 0;
      _tmp_1836 <= 0;
      _tmp_1837 <= 0;
      _tmp_1838 <= 0;
      _tmp_1839 <= 0;
      _tmp_1840 <= 0;
      _tmp_1841 <= 0;
      _tmp_1842 <= 0;
      _tmp_1843 <= 0;
      _tmp_1844 <= 0;
      _tmp_1845 <= 0;
      _tmp_1846 <= 0;
      _tmp_1847 <= 0;
      _tmp_1848 <= 0;
      _tmp_1849 <= 0;
      _tmp_1850 <= 0;
      _tmp_1851 <= 0;
      _tmp_1852 <= 0;
      _tmp_1853 <= 0;
      _tmp_1854 <= 0;
      _tmp_1855 <= 0;
      _tmp_1856 <= 0;
      _tmp_1857 <= 0;
      _tmp_1858 <= 0;
      _tmp_1859 <= 0;
      _acc_1_busy_reg <= 0;
    end else begin
      if(_acc_1_stream_oready) begin
        _acc_1_x_source_ram_renable <= 0;
        _acc_1_x_source_fifo_deq <= 0;
      end 
      _acc_1_x_idle <= _acc_1_x_idle;
      if(_acc_1_stream_oready) begin
        _acc_1_rshift_source_ram_renable <= 0;
        _acc_1_rshift_source_fifo_deq <= 0;
      end 
      _acc_1_rshift_idle <= _acc_1_rshift_idle;
      if(_acc_1_stream_oready) begin
        _acc_1_sum_sink_wenable <= 0;
        _acc_1_sum_sink_fifo_enq <= 0;
      end 
      if(_acc_1_stream_oready) begin
        _acc_1_valid_sink_wenable <= 0;
        _acc_1_valid_sink_fifo_enq <= 0;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_1 <= _acc_1_stream_ivalid;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_2 <= __acc_1_stream_ivalid_1;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_3 <= __acc_1_stream_ivalid_2;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_4 <= __acc_1_stream_ivalid_3;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_5 <= __acc_1_stream_ivalid_4;
      end 
      if(_acc_1_stream_oready) begin
        _greaterthan_data_25 <= acc_1_rshift_data > 1'sd0;
      end 
      if(_acc_1_stream_oready) begin
        _minus_data_27 <= acc_1_rshift_data - 2'sd1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready && _reduceadd_reset_cond_38) begin
        _reduceadd_data_38 <= 1'sd0;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _reduceadd_count_38 <= (_reduceadd_current_count_38 >= acc_1_size_data - 1)? 0 : _reduceadd_current_count_38 + 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _reduceadd_prev_count_max_38 <= _reduceadd_current_count_38 >= acc_1_size_data - 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _reduceadd_data_38 <= _reduceadd_current_data_38 + acc_1_x_data;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready && _pulse_reset_cond_40) begin
        _pulse_data_40 <= 1'sd0;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _pulse_count_40 <= (_pulse_current_count_40 >= acc_1_size_data - 1)? 0 : _pulse_current_count_40 + 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _pulse_prev_count_max_40 <= _pulse_current_count_40 >= acc_1_size_data - 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _pulse_data_40 <= _pulse_current_count_40 >= acc_1_size_data - 1;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_1223__variable_23 <= acc_1_rshift_data;
      end 
      if(_acc_1_stream_oready) begin
        _sll_data_29 <= 2'sd1 << _minus_data_27;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_1220_greaterthan_25 <= _greaterthan_data_25;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_1221_reduceadd_38 <= _reduceadd_data_38;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_1224__delay_1223__variable_23 <= __delay_data_1223__variable_23;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_1227_pulse_40 <= _pulse_data_40;
      end 
      if(_acc_1_stream_oready) begin
        _cond_data_35 <= (__delay_data_1220_greaterthan_25)? _sll_data_29 : 1'sd0;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_1222__delay_1221_reduceadd_38 <= __delay_data_1221_reduceadd_38;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_1225__delay_1224__delay_1223__variable_23 <= __delay_data_1224__delay_1223__variable_23;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_1228__delay_1227_pulse_40 <= __delay_data_1227_pulse_40;
      end 
      if(_acc_1_stream_oready) begin
        _plus_data_42 <= __delay_data_1222__delay_1221_reduceadd_38 + _cond_data_35;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_1226__delay_1225__delay_1224____variable_23 <= __delay_data_1225__delay_1224__delay_1223__variable_23;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_1229__delay_1228__delay_1227_pulse_40 <= __delay_data_1228__delay_1227_pulse_40;
      end 
      if(_acc_1_stream_oready) begin
        _sra_data_43 <= _plus_data_42 >>> __delay_data_1226__delay_1225__delay_1224____variable_23;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_1230__delay_1229__delay_1228__delay_1227_pulse_40 <= __delay_data_1229__delay_1228__delay_1227_pulse_40;
      end 
      if(__stream_matmul_33_stream_ivalid_14 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_37 <= __delay_data_1536__delay_1535__delay_1534____variable_1057;
      end 
      if(__stream_matmul_33_stream_ivalid_14 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_22 <= __substreamoutput_data_1218;
      end 
      if(__stream_matmul_33_stream_ivalid_14 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_23 <= __delay_data_1586__delay_1585__delay_1584___plus_1231;
      end 
      if(__stream_matmul_33_stream_ivalid_14 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_24 <= __delay_data_1563__delay_1562__delay_1561____variable_1052;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1828 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1829 <= _tmp_1828;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1830 <= _tmp_1829;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1831 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1832 <= _tmp_1831;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1833 <= _tmp_1832;
      end 
      if(_acc_1_stream_oready && _tmp_1833) begin
        __variable_wdata_37 <= 1;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1834 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1835 <= _tmp_1834;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1836 <= _tmp_1835;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1837 <= _tmp_1836;
      end 
      if(_acc_1_stream_oready && _tmp_1837) begin
        __variable_wdata_37 <= 0;
      end 
      if(_acc_1_stream_oready && 1'd0) begin
        __variable_wdata_37 <= 1;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1838 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1839 <= _tmp_1838;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1840 <= _tmp_1839;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1841 <= _tmp_1840;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1842 <= _tmp_1841;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1843 <= _tmp_1842;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1844 <= _tmp_1843;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1845 <= _acc_1_source_stop;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1846 <= _tmp_1845;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1847 <= _tmp_1846;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1848 <= _tmp_1847;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1849 <= _tmp_1848;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1850 <= _tmp_1849;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1851 <= _tmp_1850;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1852 <= _acc_1_source_busy;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1853 <= _tmp_1852;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1854 <= _tmp_1853;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1855 <= _tmp_1854;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1856 <= _tmp_1855;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1857 <= _tmp_1856;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1858 <= _tmp_1857;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1859 <= _acc_1_sink_busy;
      end 
      if(!_acc_1_sink_busy && _tmp_1859) begin
        _acc_1_busy_reg <= 0;
      end 
      if(_acc_1_source_busy) begin
        _acc_1_busy_reg <= 1;
      end 
    end
  end

  localparam _acc_1_fsm_1 = 1;
  localparam _acc_1_fsm_2 = 2;
  localparam _acc_1_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _acc_1_fsm <= _acc_1_fsm_init;
      _acc_1_source_start <= 0;
      _acc_1_source_busy <= 0;
      _acc_1_stream_ivalid <= 0;
    end else begin
      if(__stream_matmul_33_stream_ivalid_14 && _stream_matmul_33_stream_oready) begin
        _acc_1_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_busy) begin
        _acc_1_source_busy <= _stream_matmul_33_source_busy;
      end 
      if(_acc_1_stream_oready && _tmp_1830) begin
        _acc_1_stream_ivalid <= 1;
      end 
      if(_acc_1_stream_oready && 1'd0) begin
        _acc_1_stream_ivalid <= 0;
      end 
      case(_acc_1_fsm)
        _acc_1_fsm_init: begin
          if(_acc_1_run_flag) begin
            _acc_1_source_start <= 1;
          end 
          if(_acc_1_run_flag) begin
            _acc_1_fsm <= _acc_1_fsm_1;
          end 
        end
        _acc_1_fsm_1: begin
          if(_acc_1_source_start && _acc_1_stream_oready) begin
            _acc_1_source_start <= 0;
            _acc_1_source_busy <= 1;
          end 
          if(_acc_1_source_start && _acc_1_stream_oready) begin
            _acc_1_fsm <= _acc_1_fsm_2;
          end 
        end
        _acc_1_fsm_2: begin
          if(_acc_1_stream_oready) begin
            _acc_1_fsm <= _acc_1_fsm_3;
          end 
        end
        _acc_1_fsm_3: begin
          if(_acc_1_stream_oready && 1'd0) begin
            _acc_1_source_busy <= 0;
          end 
          if(_acc_1_stream_oready && 1'd0 && _acc_1_run_flag) begin
            _acc_1_source_start <= 1;
          end 
          if(_acc_1_stream_oready && 1'd0) begin
            _acc_1_fsm <= _acc_1_fsm_init;
          end 
          if(_acc_1_stream_oready && 1'd0 && _acc_1_run_flag) begin
            _acc_1_fsm <= _acc_1_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_2_var0_source_ram_renable <= 0;
      _add_tree_2_var0_source_fifo_deq <= 0;
      _add_tree_2_var0_idle <= 1;
      _add_tree_2_sum_sink_wenable <= 0;
      _add_tree_2_sum_sink_fifo_enq <= 0;
      __variable_wdata_44 <= 0;
      _tmp_1509 <= 0;
      _tmp_1510 <= 0;
      _tmp_1511 <= 0;
      _tmp_1512 <= 0;
      _tmp_1513 <= 0;
      _tmp_1514 <= 0;
      _tmp_1515 <= 0;
      _tmp_1516 <= 0;
      _tmp_1517 <= 0;
      _tmp_1518 <= 0;
      _add_tree_2_busy_reg <= 0;
    end else begin
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_var0_source_ram_renable <= 0;
        _add_tree_2_var0_source_fifo_deq <= 0;
      end 
      _add_tree_2_var0_idle <= _add_tree_2_var0_idle;
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_sum_sink_wenable <= 0;
        _add_tree_2_sum_sink_fifo_enq <= 0;
      end 
      if(__stream_matmul_23_stream_ivalid_10 && _stream_matmul_23_stream_oready) begin
        __variable_wdata_44 <= __substreamoutput_data_1036;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1509 <= _add_tree_2_source_start;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1510 <= _tmp_1509;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1511 <= _tmp_1510;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1512 <= _add_tree_2_source_start;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1513 <= _tmp_1512;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1514 <= _add_tree_2_source_stop;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1515 <= _tmp_1514;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1516 <= _add_tree_2_source_busy;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1517 <= _tmp_1516;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1518 <= _add_tree_2_sink_busy;
      end 
      if(!_add_tree_2_sink_busy && _tmp_1518) begin
        _add_tree_2_busy_reg <= 0;
      end 
      if(_add_tree_2_source_busy) begin
        _add_tree_2_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_2_fsm_1 = 1;
  localparam _add_tree_2_fsm_2 = 2;
  localparam _add_tree_2_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_2_fsm <= _add_tree_2_fsm_init;
      _add_tree_2_source_start <= 0;
      _add_tree_2_source_busy <= 0;
      _add_tree_2_stream_ivalid <= 0;
    end else begin
      if(__stream_matmul_23_stream_ivalid_10 && _stream_matmul_23_stream_oready) begin
        _add_tree_2_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_23_stream_oready && _stream_matmul_23_busy) begin
        _add_tree_2_source_busy <= _stream_matmul_23_source_busy;
      end 
      if(_add_tree_2_stream_oready && _tmp_1511) begin
        _add_tree_2_stream_ivalid <= 1;
      end 
      if(_add_tree_2_stream_oready && 1'd0) begin
        _add_tree_2_stream_ivalid <= 0;
      end 
      case(_add_tree_2_fsm)
        _add_tree_2_fsm_init: begin
          if(_add_tree_2_run_flag) begin
            _add_tree_2_source_start <= 1;
          end 
          if(_add_tree_2_run_flag) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_1;
          end 
        end
        _add_tree_2_fsm_1: begin
          if(_add_tree_2_source_start && _add_tree_2_stream_oready) begin
            _add_tree_2_source_start <= 0;
            _add_tree_2_source_busy <= 1;
          end 
          if(_add_tree_2_source_start && _add_tree_2_stream_oready) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_2;
          end 
        end
        _add_tree_2_fsm_2: begin
          if(_add_tree_2_stream_oready) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_3;
          end 
        end
        _add_tree_2_fsm_3: begin
          if(_add_tree_2_stream_oready && 1'd0) begin
            _add_tree_2_source_busy <= 0;
          end 
          if(_add_tree_2_stream_oready && 1'd0 && _add_tree_2_run_flag) begin
            _add_tree_2_source_start <= 1;
          end 
          if(_add_tree_2_stream_oready && 1'd0) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_init;
          end 
          if(_add_tree_2_stream_oready && 1'd0 && _add_tree_2_run_flag) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_3_var0_source_ram_renable <= 0;
      _add_tree_3_var0_source_fifo_deq <= 0;
      _add_tree_3_var0_idle <= 1;
      _add_tree_3_var1_source_ram_renable <= 0;
      _add_tree_3_var1_source_fifo_deq <= 0;
      _add_tree_3_var1_idle <= 1;
      _add_tree_3_sum_sink_wenable <= 0;
      _add_tree_3_sum_sink_fifo_enq <= 0;
      __add_tree_3_stream_ivalid_1 <= 0;
      __plusn_data_49 <= 0;
      __variable_wdata_46 <= 0;
      __variable_wdata_47 <= 0;
      _tmp_1802 <= 0;
      _tmp_1803 <= 0;
      _tmp_1804 <= 0;
      _tmp_1805 <= 0;
      _tmp_1806 <= 0;
      _tmp_1807 <= 0;
      _tmp_1808 <= 0;
      _tmp_1809 <= 0;
      _tmp_1810 <= 0;
      _tmp_1811 <= 0;
      _tmp_1812 <= 0;
      _tmp_1813 <= 0;
      _tmp_1814 <= 0;
      _add_tree_3_busy_reg <= 0;
    end else begin
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_var0_source_ram_renable <= 0;
        _add_tree_3_var0_source_fifo_deq <= 0;
      end 
      _add_tree_3_var0_idle <= _add_tree_3_var0_idle;
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_var1_source_ram_renable <= 0;
        _add_tree_3_var1_source_fifo_deq <= 0;
      end 
      _add_tree_3_var1_idle <= _add_tree_3_var1_idle;
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_sum_sink_wenable <= 0;
        _add_tree_3_sum_sink_fifo_enq <= 0;
      end 
      if(_add_tree_3_stream_oready) begin
        __add_tree_3_stream_ivalid_1 <= _add_tree_3_stream_ivalid;
      end 
      if(_add_tree_3_stream_oready) begin
        __plusn_data_49 <= add_tree_3_var0_data + add_tree_3_var1_data + 1'sd0;
      end 
      if(__stream_matmul_33_stream_ivalid_12 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_46 <= __substreamoutput_data_1190;
      end 
      if(__stream_matmul_33_stream_ivalid_12 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_47 <= __substreamoutput_data_1195;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1802 <= _add_tree_3_source_start;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1803 <= _tmp_1802;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1804 <= _tmp_1803;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1805 <= _add_tree_3_source_start;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1806 <= _tmp_1805;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1807 <= _tmp_1806;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1808 <= _add_tree_3_source_stop;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1809 <= _tmp_1808;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1810 <= _tmp_1809;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1811 <= _add_tree_3_source_busy;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1812 <= _tmp_1811;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1813 <= _tmp_1812;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1814 <= _add_tree_3_sink_busy;
      end 
      if(!_add_tree_3_sink_busy && _tmp_1814) begin
        _add_tree_3_busy_reg <= 0;
      end 
      if(_add_tree_3_source_busy) begin
        _add_tree_3_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_3_fsm_1 = 1;
  localparam _add_tree_3_fsm_2 = 2;
  localparam _add_tree_3_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_3_fsm <= _add_tree_3_fsm_init;
      _add_tree_3_source_start <= 0;
      _add_tree_3_source_busy <= 0;
      _add_tree_3_stream_ivalid <= 0;
    end else begin
      if(__stream_matmul_33_stream_ivalid_12 && _stream_matmul_33_stream_oready) begin
        _add_tree_3_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_busy) begin
        _add_tree_3_source_busy <= _stream_matmul_33_source_busy;
      end 
      if(_add_tree_3_stream_oready && _tmp_1804) begin
        _add_tree_3_stream_ivalid <= 1;
      end 
      if(_add_tree_3_stream_oready && 1'd0) begin
        _add_tree_3_stream_ivalid <= 0;
      end 
      case(_add_tree_3_fsm)
        _add_tree_3_fsm_init: begin
          if(_add_tree_3_run_flag) begin
            _add_tree_3_source_start <= 1;
          end 
          if(_add_tree_3_run_flag) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_1;
          end 
        end
        _add_tree_3_fsm_1: begin
          if(_add_tree_3_source_start && _add_tree_3_stream_oready) begin
            _add_tree_3_source_start <= 0;
            _add_tree_3_source_busy <= 1;
          end 
          if(_add_tree_3_source_start && _add_tree_3_stream_oready) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_2;
          end 
        end
        _add_tree_3_fsm_2: begin
          if(_add_tree_3_stream_oready) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_3;
          end 
        end
        _add_tree_3_fsm_3: begin
          if(_add_tree_3_stream_oready && 1'd0) begin
            _add_tree_3_source_busy <= 0;
          end 
          if(_add_tree_3_stream_oready && 1'd0 && _add_tree_3_run_flag) begin
            _add_tree_3_source_start <= 1;
          end 
          if(_add_tree_3_stream_oready && 1'd0) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_init;
          end 
          if(_add_tree_3_stream_oready && 1'd0 && _add_tree_3_run_flag) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_4_var0_source_ram_renable <= 0;
      _add_tree_4_var0_source_fifo_deq <= 0;
      _add_tree_4_var0_idle <= 1;
      _add_tree_4_var1_source_ram_renable <= 0;
      _add_tree_4_var1_source_fifo_deq <= 0;
      _add_tree_4_var1_idle <= 1;
      _add_tree_4_sum_sink_wenable <= 0;
      _add_tree_4_sum_sink_fifo_enq <= 0;
      __add_tree_4_stream_ivalid_1 <= 0;
      __plusn_data_53 <= 0;
      __variable_wdata_50 <= 0;
      __variable_wdata_51 <= 0;
      _tmp_1815 <= 0;
      _tmp_1816 <= 0;
      _tmp_1817 <= 0;
      _tmp_1818 <= 0;
      _tmp_1819 <= 0;
      _tmp_1820 <= 0;
      _tmp_1821 <= 0;
      _tmp_1822 <= 0;
      _tmp_1823 <= 0;
      _tmp_1824 <= 0;
      _tmp_1825 <= 0;
      _tmp_1826 <= 0;
      _tmp_1827 <= 0;
      _add_tree_4_busy_reg <= 0;
    end else begin
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var0_source_ram_renable <= 0;
        _add_tree_4_var0_source_fifo_deq <= 0;
      end 
      _add_tree_4_var0_idle <= _add_tree_4_var0_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var1_source_ram_renable <= 0;
        _add_tree_4_var1_source_fifo_deq <= 0;
      end 
      _add_tree_4_var1_idle <= _add_tree_4_var1_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_sum_sink_wenable <= 0;
        _add_tree_4_sum_sink_fifo_enq <= 0;
      end 
      if(_add_tree_4_stream_oready) begin
        __add_tree_4_stream_ivalid_1 <= _add_tree_4_stream_ivalid;
      end 
      if(_add_tree_4_stream_oready) begin
        __plusn_data_53 <= add_tree_4_var0_data + add_tree_4_var1_data + 1'sd0;
      end 
      if(__stream_matmul_33_stream_ivalid_12 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_50 <= __substreamoutput_data_1211;
      end 
      if(__stream_matmul_33_stream_ivalid_12 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_51 <= __substreamoutput_data_1216;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1815 <= _add_tree_4_source_start;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1816 <= _tmp_1815;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1817 <= _tmp_1816;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1818 <= _add_tree_4_source_start;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1819 <= _tmp_1818;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1820 <= _tmp_1819;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1821 <= _add_tree_4_source_stop;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1822 <= _tmp_1821;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1823 <= _tmp_1822;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1824 <= _add_tree_4_source_busy;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1825 <= _tmp_1824;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1826 <= _tmp_1825;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1827 <= _add_tree_4_sink_busy;
      end 
      if(!_add_tree_4_sink_busy && _tmp_1827) begin
        _add_tree_4_busy_reg <= 0;
      end 
      if(_add_tree_4_source_busy) begin
        _add_tree_4_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_4_fsm_1 = 1;
  localparam _add_tree_4_fsm_2 = 2;
  localparam _add_tree_4_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_4_fsm <= _add_tree_4_fsm_init;
      _add_tree_4_source_start <= 0;
      _add_tree_4_source_busy <= 0;
      _add_tree_4_stream_ivalid <= 0;
    end else begin
      if(__stream_matmul_33_stream_ivalid_12 && _stream_matmul_33_stream_oready) begin
        _add_tree_4_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_busy) begin
        _add_tree_4_source_busy <= _stream_matmul_33_source_busy;
      end 
      if(_add_tree_4_stream_oready && _tmp_1817) begin
        _add_tree_4_stream_ivalid <= 1;
      end 
      if(_add_tree_4_stream_oready && 1'd0) begin
        _add_tree_4_stream_ivalid <= 0;
      end 
      case(_add_tree_4_fsm)
        _add_tree_4_fsm_init: begin
          if(_add_tree_4_run_flag) begin
            _add_tree_4_source_start <= 1;
          end 
          if(_add_tree_4_run_flag) begin
            _add_tree_4_fsm <= _add_tree_4_fsm_1;
          end 
        end
        _add_tree_4_fsm_1: begin
          if(_add_tree_4_source_start && _add_tree_4_stream_oready) begin
            _add_tree_4_source_start <= 0;
            _add_tree_4_source_busy <= 1;
          end 
          if(_add_tree_4_source_start && _add_tree_4_stream_oready) begin
            _add_tree_4_fsm <= _add_tree_4_fsm_2;
          end 
        end
        _add_tree_4_fsm_2: begin
          if(_add_tree_4_stream_oready) begin
            _add_tree_4_fsm <= _add_tree_4_fsm_3;
          end 
        end
        _add_tree_4_fsm_3: begin
          if(_add_tree_4_stream_oready && 1'd0) begin
            _add_tree_4_source_busy <= 0;
          end 
          if(_add_tree_4_stream_oready && 1'd0 && _add_tree_4_run_flag) begin
            _add_tree_4_source_start <= 1;
          end 
          if(_add_tree_4_stream_oready && 1'd0) begin
            _add_tree_4_fsm <= _add_tree_4_fsm_init;
          end 
          if(_add_tree_4_stream_oready && 1'd0 && _add_tree_4_run_flag) begin
            _add_tree_4_fsm <= _add_tree_4_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_5_var0_source_ram_renable <= 0;
      _add_tree_5_var0_source_fifo_deq <= 0;
      _add_tree_5_var0_idle <= 1;
      _add_tree_5_var1_source_ram_renable <= 0;
      _add_tree_5_var1_source_fifo_deq <= 0;
      _add_tree_5_var1_idle <= 1;
      _add_tree_5_var2_source_ram_renable <= 0;
      _add_tree_5_var2_source_fifo_deq <= 0;
      _add_tree_5_var2_idle <= 1;
      _add_tree_5_var3_source_ram_renable <= 0;
      _add_tree_5_var3_source_fifo_deq <= 0;
      _add_tree_5_var3_idle <= 1;
      _add_tree_5_var4_source_ram_renable <= 0;
      _add_tree_5_var4_source_fifo_deq <= 0;
      _add_tree_5_var4_idle <= 1;
      _add_tree_5_var5_source_ram_renable <= 0;
      _add_tree_5_var5_source_fifo_deq <= 0;
      _add_tree_5_var5_idle <= 1;
      _add_tree_5_var6_source_ram_renable <= 0;
      _add_tree_5_var6_source_fifo_deq <= 0;
      _add_tree_5_var6_idle <= 1;
      _add_tree_5_var7_source_ram_renable <= 0;
      _add_tree_5_var7_source_fifo_deq <= 0;
      _add_tree_5_var7_idle <= 1;
      _add_tree_5_var8_source_ram_renable <= 0;
      _add_tree_5_var8_source_fifo_deq <= 0;
      _add_tree_5_var8_idle <= 1;
      _add_tree_5_sum_sink_wenable <= 0;
      _add_tree_5_sum_sink_fifo_enq <= 0;
      __add_tree_5_stream_ivalid_1 <= 0;
      __add_tree_5_stream_ivalid_2 <= 0;
      __plusn_data_64 <= 0;
      __plusn_data_65 <= 0;
      __plusn_data_66 <= 0;
      __plusn_data_67 <= 0;
      __variable_wdata_54 <= 0;
      __variable_wdata_55 <= 0;
      __variable_wdata_56 <= 0;
      __variable_wdata_57 <= 0;
      __variable_wdata_58 <= 0;
      __variable_wdata_59 <= 0;
      __variable_wdata_60 <= 0;
      __variable_wdata_61 <= 0;
      __variable_wdata_62 <= 0;
      _tmp_935 <= 0;
      _tmp_936 <= 0;
      _tmp_937 <= 0;
      _tmp_938 <= 0;
      _tmp_939 <= 0;
      _tmp_940 <= 0;
      _tmp_941 <= 0;
      _tmp_942 <= 0;
      _tmp_943 <= 0;
      _tmp_944 <= 0;
      _tmp_945 <= 0;
      _tmp_946 <= 0;
      _tmp_947 <= 0;
      _tmp_948 <= 0;
      _tmp_949 <= 0;
      _tmp_950 <= 0;
      _add_tree_5_busy_reg <= 0;
    end else begin
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var0_source_ram_renable <= 0;
        _add_tree_5_var0_source_fifo_deq <= 0;
      end 
      _add_tree_5_var0_idle <= _add_tree_5_var0_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var1_source_ram_renable <= 0;
        _add_tree_5_var1_source_fifo_deq <= 0;
      end 
      _add_tree_5_var1_idle <= _add_tree_5_var1_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var2_source_ram_renable <= 0;
        _add_tree_5_var2_source_fifo_deq <= 0;
      end 
      _add_tree_5_var2_idle <= _add_tree_5_var2_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var3_source_ram_renable <= 0;
        _add_tree_5_var3_source_fifo_deq <= 0;
      end 
      _add_tree_5_var3_idle <= _add_tree_5_var3_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var4_source_ram_renable <= 0;
        _add_tree_5_var4_source_fifo_deq <= 0;
      end 
      _add_tree_5_var4_idle <= _add_tree_5_var4_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var5_source_ram_renable <= 0;
        _add_tree_5_var5_source_fifo_deq <= 0;
      end 
      _add_tree_5_var5_idle <= _add_tree_5_var5_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var6_source_ram_renable <= 0;
        _add_tree_5_var6_source_fifo_deq <= 0;
      end 
      _add_tree_5_var6_idle <= _add_tree_5_var6_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var7_source_ram_renable <= 0;
        _add_tree_5_var7_source_fifo_deq <= 0;
      end 
      _add_tree_5_var7_idle <= _add_tree_5_var7_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var8_source_ram_renable <= 0;
        _add_tree_5_var8_source_fifo_deq <= 0;
      end 
      _add_tree_5_var8_idle <= _add_tree_5_var8_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_sum_sink_wenable <= 0;
        _add_tree_5_sum_sink_fifo_enq <= 0;
      end 
      if(_add_tree_5_stream_oready) begin
        __add_tree_5_stream_ivalid_1 <= _add_tree_5_stream_ivalid;
      end 
      if(_add_tree_5_stream_oready) begin
        __add_tree_5_stream_ivalid_2 <= __add_tree_5_stream_ivalid_1;
      end 
      if(_add_tree_5_stream_oready) begin
        __plusn_data_64 <= add_tree_5_var0_data + add_tree_5_var1_data + add_tree_5_var2_data;
      end 
      if(_add_tree_5_stream_oready) begin
        __plusn_data_65 <= add_tree_5_var3_data + add_tree_5_var4_data + add_tree_5_var5_data;
      end 
      if(_add_tree_5_stream_oready) begin
        __plusn_data_66 <= add_tree_5_var6_data + add_tree_5_var7_data + add_tree_5_var8_data;
      end 
      if(_add_tree_5_stream_oready) begin
        __plusn_data_67 <= __plusn_data_64 + __plusn_data_65 + __plusn_data_66;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_54 <= __substreamoutput_data_735;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_55 <= __substreamoutput_data_754;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_56 <= __substreamoutput_data_773;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_57 <= __substreamoutput_data_792;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_58 <= __substreamoutput_data_811;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_59 <= __substreamoutput_data_830;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_60 <= __substreamoutput_data_849;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_61 <= __substreamoutput_data_868;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_62 <= __substreamoutput_data_887;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_935 <= _add_tree_5_source_start;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_936 <= _tmp_935;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_937 <= _tmp_936;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_938 <= _add_tree_5_source_start;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_939 <= _tmp_938;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_940 <= _tmp_939;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_941 <= _tmp_940;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_942 <= _add_tree_5_source_stop;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_943 <= _tmp_942;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_944 <= _tmp_943;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_945 <= _tmp_944;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_946 <= _add_tree_5_source_busy;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_947 <= _tmp_946;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_948 <= _tmp_947;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_949 <= _tmp_948;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_950 <= _add_tree_5_sink_busy;
      end 
      if(!_add_tree_5_sink_busy && _tmp_950) begin
        _add_tree_5_busy_reg <= 0;
      end 
      if(_add_tree_5_source_busy) begin
        _add_tree_5_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_5_fsm_1 = 1;
  localparam _add_tree_5_fsm_2 = 2;
  localparam _add_tree_5_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_5_fsm <= _add_tree_5_fsm_init;
      _add_tree_5_source_start <= 0;
      _add_tree_5_source_busy <= 0;
      _add_tree_5_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        _add_tree_5_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _add_tree_5_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_add_tree_5_stream_oready && _tmp_937) begin
        _add_tree_5_stream_ivalid <= 1;
      end 
      if(_add_tree_5_stream_oready && 1'd0) begin
        _add_tree_5_stream_ivalid <= 0;
      end 
      case(_add_tree_5_fsm)
        _add_tree_5_fsm_init: begin
          if(_add_tree_5_run_flag) begin
            _add_tree_5_source_start <= 1;
          end 
          if(_add_tree_5_run_flag) begin
            _add_tree_5_fsm <= _add_tree_5_fsm_1;
          end 
        end
        _add_tree_5_fsm_1: begin
          if(_add_tree_5_source_start && _add_tree_5_stream_oready) begin
            _add_tree_5_source_start <= 0;
            _add_tree_5_source_busy <= 1;
          end 
          if(_add_tree_5_source_start && _add_tree_5_stream_oready) begin
            _add_tree_5_fsm <= _add_tree_5_fsm_2;
          end 
        end
        _add_tree_5_fsm_2: begin
          if(_add_tree_5_stream_oready) begin
            _add_tree_5_fsm <= _add_tree_5_fsm_3;
          end 
        end
        _add_tree_5_fsm_3: begin
          if(_add_tree_5_stream_oready && 1'd0) begin
            _add_tree_5_source_busy <= 0;
          end 
          if(_add_tree_5_stream_oready && 1'd0 && _add_tree_5_run_flag) begin
            _add_tree_5_source_start <= 1;
          end 
          if(_add_tree_5_stream_oready && 1'd0) begin
            _add_tree_5_fsm <= _add_tree_5_fsm_init;
          end 
          if(_add_tree_5_stream_oready && 1'd0 && _add_tree_5_run_flag) begin
            _add_tree_5_fsm <= _add_tree_5_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_6_x_source_ram_renable <= 0;
      _mul_rshift_round_clip_6_x_source_fifo_deq <= 0;
      _mul_rshift_round_clip_6_x_idle <= 1;
      _mul_rshift_round_clip_6_y_source_ram_renable <= 0;
      _mul_rshift_round_clip_6_y_source_fifo_deq <= 0;
      _mul_rshift_round_clip_6_y_idle <= 1;
      _mul_rshift_round_clip_6_rshift_source_ram_renable <= 0;
      _mul_rshift_round_clip_6_rshift_source_fifo_deq <= 0;
      _mul_rshift_round_clip_6_rshift_idle <= 1;
      _mul_rshift_round_clip_6_z_sink_wenable <= 0;
      _mul_rshift_round_clip_6_z_sink_fifo_enq <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_1 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_2 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_3 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_4 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_5 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_6 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_7 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_8 <= 0;
      _times_mul_odata_reg_71 <= 0;
      __delay_data_907_sll_77 <= 0;
      __delay_data_911__variable_70 <= 0;
      __delay_data_915_eq_89 <= 0;
      __delay_data_908__delay_907_sll_77 <= 0;
      __delay_data_912__delay_911__variable_70 <= 0;
      __delay_data_916__delay_915_eq_89 <= 0;
      __delay_data_909__delay_908__delay_907_sll_77 <= 0;
      __delay_data_913__delay_912__delay_911__variable_70 <= 0;
      __delay_data_917__delay_916__delay_915_eq_89 <= 0;
      __delay_data_910__delay_909__delay_908__delay_907_sll_77 <= 0;
      __delay_data_914__delay_913__delay_912__delay_911__variable_70 <= 0;
      __delay_data_918__delay_917__delay_916__delay_915_eq_89 <= 0;
      _cond_data_90 <= 0;
      _greaterthan_data_91 <= 0;
      _lessthan_data_95 <= 0;
      _greatereq_data_99 <= 0;
      __delay_data_919_cond_90 <= 0;
      _cond_data_93 <= 0;
      _cond_data_97 <= 0;
      __delay_data_920_greatereq_99 <= 0;
      _cond_data_101 <= 0;
      __variable_wdata_68 <= 0;
      __variable_wdata_69 <= 0;
      __variable_wdata_70 <= 0;
      _tmp_983 <= 0;
      _tmp_984 <= 0;
      _tmp_985 <= 0;
      _tmp_986 <= 0;
      _tmp_987 <= 0;
      _tmp_988 <= 0;
      _tmp_989 <= 0;
      _tmp_990 <= 0;
      _tmp_991 <= 0;
      _tmp_992 <= 0;
      _tmp_993 <= 0;
      _tmp_994 <= 0;
      _tmp_995 <= 0;
      _tmp_996 <= 0;
      _tmp_997 <= 0;
      _tmp_998 <= 0;
      _tmp_999 <= 0;
      _tmp_1000 <= 0;
      _tmp_1001 <= 0;
      _tmp_1002 <= 0;
      _tmp_1003 <= 0;
      _tmp_1004 <= 0;
      _tmp_1005 <= 0;
      _tmp_1006 <= 0;
      _tmp_1007 <= 0;
      _tmp_1008 <= 0;
      _tmp_1009 <= 0;
      _tmp_1010 <= 0;
      _tmp_1011 <= 0;
      _tmp_1012 <= 0;
      _tmp_1013 <= 0;
      _tmp_1014 <= 0;
      _tmp_1015 <= 0;
      _tmp_1016 <= 0;
      _mul_rshift_round_clip_6_busy_reg <= 0;
    end else begin
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _mul_rshift_round_clip_6_x_source_ram_renable <= 0;
        _mul_rshift_round_clip_6_x_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_6_x_idle <= _mul_rshift_round_clip_6_x_idle;
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _mul_rshift_round_clip_6_y_source_ram_renable <= 0;
        _mul_rshift_round_clip_6_y_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_6_y_idle <= _mul_rshift_round_clip_6_y_idle;
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _mul_rshift_round_clip_6_rshift_source_ram_renable <= 0;
        _mul_rshift_round_clip_6_rshift_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_6_rshift_idle <= _mul_rshift_round_clip_6_rshift_idle;
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _mul_rshift_round_clip_6_z_sink_wenable <= 0;
        _mul_rshift_round_clip_6_z_sink_fifo_enq <= 0;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_1 <= _mul_rshift_round_clip_6_stream_ivalid;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_2 <= __mul_rshift_round_clip_6_stream_ivalid_1;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_3 <= __mul_rshift_round_clip_6_stream_ivalid_2;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_4 <= __mul_rshift_round_clip_6_stream_ivalid_3;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_5 <= __mul_rshift_round_clip_6_stream_ivalid_4;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_6 <= __mul_rshift_round_clip_6_stream_ivalid_5;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_7 <= __mul_rshift_round_clip_6_stream_ivalid_6;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_8 <= __mul_rshift_round_clip_6_stream_ivalid_7;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _times_mul_odata_reg_71 <= _times_mul_odata_71;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_907_sll_77 <= _sll_data_77;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_911__variable_70 <= mul_rshift_round_clip_6_rshift_data;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_915_eq_89 <= _eq_data_89;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_908__delay_907_sll_77 <= __delay_data_907_sll_77;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_912__delay_911__variable_70 <= __delay_data_911__variable_70;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_916__delay_915_eq_89 <= __delay_data_915_eq_89;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_909__delay_908__delay_907_sll_77 <= __delay_data_908__delay_907_sll_77;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_913__delay_912__delay_911__variable_70 <= __delay_data_912__delay_911__variable_70;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_917__delay_916__delay_915_eq_89 <= __delay_data_916__delay_915_eq_89;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_910__delay_909__delay_908__delay_907_sll_77 <= __delay_data_909__delay_908__delay_907_sll_77;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_914__delay_913__delay_912__delay_911__variable_70 <= __delay_data_913__delay_912__delay_911__variable_70;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_918__delay_917__delay_916__delay_915_eq_89 <= __delay_data_917__delay_916__delay_915_eq_89;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _cond_data_90 <= (__delay_data_918__delay_917__delay_916__delay_915_eq_89)? _times_data_71 : _sra_data_87;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _greaterthan_data_91 <= _cond_data_90 > 16'sd32767;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _lessthan_data_95 <= _cond_data_90 < -16'sd32767;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _greatereq_data_99 <= _cond_data_90 >= 1'sd0;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_919_cond_90 <= _cond_data_90;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _cond_data_93 <= (_greaterthan_data_91)? 16'sd32767 : __delay_data_919_cond_90;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _cond_data_97 <= (_lessthan_data_95)? -16'sd32767 : __delay_data_919_cond_90;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_920_greatereq_99 <= _greatereq_data_99;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _cond_data_101 <= (__delay_data_920_greatereq_99)? _cond_data_93 : _cond_data_97;
      end 
      if(__stream_conv2d_4_stream_ivalid_20 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_68 <= _plus_data_905;
      end 
      if(__stream_conv2d_4_stream_ivalid_20 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_69 <= __delay_data_1357__delay_1356__delay_1355__delay_1354___cond_367;
      end 
      if(__stream_conv2d_4_stream_ivalid_20 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_70 <= __delay_data_1376__delay_1375__delay_1374__delay_1373___plus_921;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_983 <= _mul_rshift_round_clip_6_source_start;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_984 <= _tmp_983;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_985 <= _tmp_984;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_986 <= _mul_rshift_round_clip_6_source_start;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_987 <= _tmp_986;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_988 <= _tmp_987;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_989 <= _tmp_988;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_990 <= _tmp_989;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_991 <= _tmp_990;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_992 <= _tmp_991;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_993 <= _tmp_992;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_994 <= _tmp_993;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_995 <= _tmp_994;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_996 <= _mul_rshift_round_clip_6_source_stop;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_997 <= _tmp_996;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_998 <= _tmp_997;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_999 <= _tmp_998;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1000 <= _tmp_999;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1001 <= _tmp_1000;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1002 <= _tmp_1001;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1003 <= _tmp_1002;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1004 <= _tmp_1003;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1005 <= _tmp_1004;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1006 <= _mul_rshift_round_clip_6_source_busy;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1007 <= _tmp_1006;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1008 <= _tmp_1007;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1009 <= _tmp_1008;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1010 <= _tmp_1009;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1011 <= _tmp_1010;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1012 <= _tmp_1011;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1013 <= _tmp_1012;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1014 <= _tmp_1013;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1015 <= _tmp_1014;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1016 <= _mul_rshift_round_clip_6_sink_busy;
      end 
      if(!_mul_rshift_round_clip_6_sink_busy && _tmp_1016) begin
        _mul_rshift_round_clip_6_busy_reg <= 0;
      end 
      if(_mul_rshift_round_clip_6_source_busy) begin
        _mul_rshift_round_clip_6_busy_reg <= 1;
      end 
      if(__stream_matmul_23_stream_ivalid_18 && _stream_matmul_23_stream_oready) begin
        __variable_wdata_68 <= _plus_data_1043;
      end 
      if(__stream_matmul_23_stream_ivalid_18 && _stream_matmul_23_stream_oready) begin
        __variable_wdata_69 <= __delay_data_1470__delay_1469__delay_1468__delay_1467___cond_984;
      end 
      if(__stream_matmul_23_stream_ivalid_18 && _stream_matmul_23_stream_oready) begin
        __variable_wdata_70 <= __delay_data_1487__delay_1486__delay_1485___plus_1045;
      end 
      if(__stream_matmul_33_stream_ivalid_21 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_68 <= _plus_data_1202;
      end 
      if(__stream_matmul_33_stream_ivalid_21 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_69 <= __delay_data_1688__delay_1687__delay_1686___cond_1095;
      end 
      if(__stream_matmul_33_stream_ivalid_21 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_70 <= __delay_data_1708__delay_1707__delay_1706___plus_1204;
      end 
    end
  end

  localparam _mul_rshift_round_clip_6_fsm_1 = 1;
  localparam _mul_rshift_round_clip_6_fsm_2 = 2;
  localparam _mul_rshift_round_clip_6_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_6_fsm <= _mul_rshift_round_clip_6_fsm_init;
      _mul_rshift_round_clip_6_source_start <= 0;
      _mul_rshift_round_clip_6_source_busy <= 0;
      _mul_rshift_round_clip_6_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_20 && _stream_conv2d_4_stream_oready) begin
        _mul_rshift_round_clip_6_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_rshift_round_clip_6_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_rshift_round_clip_6_stream_oready && _tmp_985) begin
        _mul_rshift_round_clip_6_stream_ivalid <= 1;
      end 
      if(_mul_rshift_round_clip_6_stream_oready && 1'd0) begin
        _mul_rshift_round_clip_6_stream_ivalid <= 0;
      end 
      if(__stream_matmul_23_stream_ivalid_18 && _stream_matmul_23_stream_oready) begin
        _mul_rshift_round_clip_6_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_23_stream_oready && _stream_matmul_23_busy) begin
        _mul_rshift_round_clip_6_source_busy <= _stream_matmul_23_source_busy;
      end 
      if(__stream_matmul_33_stream_ivalid_21 && _stream_matmul_33_stream_oready) begin
        _mul_rshift_round_clip_6_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_busy) begin
        _mul_rshift_round_clip_6_source_busy <= _stream_matmul_33_source_busy;
      end 
      case(_mul_rshift_round_clip_6_fsm)
        _mul_rshift_round_clip_6_fsm_init: begin
          if(_mul_rshift_round_clip_6_run_flag) begin
            _mul_rshift_round_clip_6_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_6_run_flag) begin
            _mul_rshift_round_clip_6_fsm <= _mul_rshift_round_clip_6_fsm_1;
          end 
        end
        _mul_rshift_round_clip_6_fsm_1: begin
          if(_mul_rshift_round_clip_6_source_start && _mul_rshift_round_clip_6_stream_oready) begin
            _mul_rshift_round_clip_6_source_start <= 0;
            _mul_rshift_round_clip_6_source_busy <= 1;
          end 
          if(_mul_rshift_round_clip_6_source_start && _mul_rshift_round_clip_6_stream_oready) begin
            _mul_rshift_round_clip_6_fsm <= _mul_rshift_round_clip_6_fsm_2;
          end 
        end
        _mul_rshift_round_clip_6_fsm_2: begin
          if(_mul_rshift_round_clip_6_stream_oready) begin
            _mul_rshift_round_clip_6_fsm <= _mul_rshift_round_clip_6_fsm_3;
          end 
        end
        _mul_rshift_round_clip_6_fsm_3: begin
          if(_mul_rshift_round_clip_6_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_6_source_busy <= 0;
          end 
          if(_mul_rshift_round_clip_6_stream_oready && 1'd0 && _mul_rshift_round_clip_6_run_flag) begin
            _mul_rshift_round_clip_6_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_6_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_6_fsm <= _mul_rshift_round_clip_6_fsm_init;
          end 
          if(_mul_rshift_round_clip_6_stream_oready && 1'd0 && _mul_rshift_round_clip_6_run_flag) begin
            _mul_rshift_round_clip_6_fsm <= _mul_rshift_round_clip_6_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_7_x_source_ram_renable <= 0;
      _mul_rshift_round_clip_7_x_source_fifo_deq <= 0;
      _mul_rshift_round_clip_7_x_idle <= 1;
      _mul_rshift_round_clip_7_y_source_ram_renable <= 0;
      _mul_rshift_round_clip_7_y_source_fifo_deq <= 0;
      _mul_rshift_round_clip_7_y_idle <= 1;
      _mul_rshift_round_clip_7_rshift_source_ram_renable <= 0;
      _mul_rshift_round_clip_7_rshift_source_fifo_deq <= 0;
      _mul_rshift_round_clip_7_rshift_idle <= 1;
      _mul_rshift_round_clip_7_z_sink_wenable <= 0;
      _mul_rshift_round_clip_7_z_sink_fifo_enq <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_1 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_2 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_3 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_4 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_5 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_6 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_7 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_8 <= 0;
      _times_mul_odata_reg_105 <= 0;
      __delay_data_1236_sll_111 <= 0;
      __delay_data_1240__variable_104 <= 0;
      __delay_data_1244_eq_123 <= 0;
      __delay_data_1237__delay_1236_sll_111 <= 0;
      __delay_data_1241__delay_1240__variable_104 <= 0;
      __delay_data_1245__delay_1244_eq_123 <= 0;
      __delay_data_1238__delay_1237__delay_1236_sll_111 <= 0;
      __delay_data_1242__delay_1241__delay_1240__variable_104 <= 0;
      __delay_data_1246__delay_1245__delay_1244_eq_123 <= 0;
      __delay_data_1239__delay_1238__delay_1237__delay_1236_sll_111 <= 0;
      __delay_data_1243__delay_1242__delay_1241____variable_104 <= 0;
      __delay_data_1247__delay_1246__delay_1245__delay_1244_eq_123 <= 0;
      _cond_data_124 <= 0;
      _greaterthan_data_125 <= 0;
      _lessthan_data_129 <= 0;
      _greatereq_data_133 <= 0;
      __delay_data_1248_cond_124 <= 0;
      _cond_data_127 <= 0;
      _cond_data_131 <= 0;
      __delay_data_1249_greatereq_133 <= 0;
      _cond_data_135 <= 0;
      __variable_wdata_102 <= 0;
      __variable_wdata_103 <= 0;
      __variable_wdata_104 <= 0;
      _tmp_1860 <= 0;
      _tmp_1861 <= 0;
      _tmp_1862 <= 0;
      _tmp_1863 <= 0;
      _tmp_1864 <= 0;
      _tmp_1865 <= 0;
      _tmp_1866 <= 0;
      _tmp_1867 <= 0;
      _tmp_1868 <= 0;
      _tmp_1869 <= 0;
      _tmp_1870 <= 0;
      _tmp_1871 <= 0;
      _tmp_1872 <= 0;
      _tmp_1873 <= 0;
      _tmp_1874 <= 0;
      _tmp_1875 <= 0;
      _tmp_1876 <= 0;
      _tmp_1877 <= 0;
      _tmp_1878 <= 0;
      _tmp_1879 <= 0;
      _tmp_1880 <= 0;
      _tmp_1881 <= 0;
      _tmp_1882 <= 0;
      _tmp_1883 <= 0;
      _tmp_1884 <= 0;
      _tmp_1885 <= 0;
      _tmp_1886 <= 0;
      _tmp_1887 <= 0;
      _tmp_1888 <= 0;
      _tmp_1889 <= 0;
      _tmp_1890 <= 0;
      _tmp_1891 <= 0;
      _tmp_1892 <= 0;
      _tmp_1893 <= 0;
      _mul_rshift_round_clip_7_busy_reg <= 0;
    end else begin
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _mul_rshift_round_clip_7_x_source_ram_renable <= 0;
        _mul_rshift_round_clip_7_x_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_7_x_idle <= _mul_rshift_round_clip_7_x_idle;
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _mul_rshift_round_clip_7_y_source_ram_renable <= 0;
        _mul_rshift_round_clip_7_y_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_7_y_idle <= _mul_rshift_round_clip_7_y_idle;
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _mul_rshift_round_clip_7_rshift_source_ram_renable <= 0;
        _mul_rshift_round_clip_7_rshift_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_7_rshift_idle <= _mul_rshift_round_clip_7_rshift_idle;
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _mul_rshift_round_clip_7_z_sink_wenable <= 0;
        _mul_rshift_round_clip_7_z_sink_fifo_enq <= 0;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_1 <= _mul_rshift_round_clip_7_stream_ivalid;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_2 <= __mul_rshift_round_clip_7_stream_ivalid_1;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_3 <= __mul_rshift_round_clip_7_stream_ivalid_2;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_4 <= __mul_rshift_round_clip_7_stream_ivalid_3;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_5 <= __mul_rshift_round_clip_7_stream_ivalid_4;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_6 <= __mul_rshift_round_clip_7_stream_ivalid_5;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_7 <= __mul_rshift_round_clip_7_stream_ivalid_6;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_8 <= __mul_rshift_round_clip_7_stream_ivalid_7;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _times_mul_odata_reg_105 <= _times_mul_odata_105;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1236_sll_111 <= _sll_data_111;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1240__variable_104 <= mul_rshift_round_clip_7_rshift_data;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1244_eq_123 <= _eq_data_123;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1237__delay_1236_sll_111 <= __delay_data_1236_sll_111;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1241__delay_1240__variable_104 <= __delay_data_1240__variable_104;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1245__delay_1244_eq_123 <= __delay_data_1244_eq_123;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1238__delay_1237__delay_1236_sll_111 <= __delay_data_1237__delay_1236_sll_111;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1242__delay_1241__delay_1240__variable_104 <= __delay_data_1241__delay_1240__variable_104;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1246__delay_1245__delay_1244_eq_123 <= __delay_data_1245__delay_1244_eq_123;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1239__delay_1238__delay_1237__delay_1236_sll_111 <= __delay_data_1238__delay_1237__delay_1236_sll_111;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1243__delay_1242__delay_1241____variable_104 <= __delay_data_1242__delay_1241__delay_1240__variable_104;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1247__delay_1246__delay_1245__delay_1244_eq_123 <= __delay_data_1246__delay_1245__delay_1244_eq_123;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _cond_data_124 <= (__delay_data_1247__delay_1246__delay_1245__delay_1244_eq_123)? _times_data_105 : _sra_data_121;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _greaterthan_data_125 <= _cond_data_124 > 16'sd32767;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _lessthan_data_129 <= _cond_data_124 < -16'sd32767;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _greatereq_data_133 <= _cond_data_124 >= 1'sd0;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1248_cond_124 <= _cond_data_124;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _cond_data_127 <= (_greaterthan_data_125)? 16'sd32767 : __delay_data_1248_cond_124;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _cond_data_131 <= (_lessthan_data_129)? -16'sd32767 : __delay_data_1248_cond_124;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_1249_greatereq_133 <= _greatereq_data_133;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _cond_data_135 <= (__delay_data_1249_greatereq_133)? _cond_data_127 : _cond_data_131;
      end 
      if(__stream_matmul_33_stream_ivalid_21 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_102 <= _plus_data_1234;
      end 
      if(__stream_matmul_33_stream_ivalid_21 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_103 <= __delay_data_1627__delay_1626__delay_1625___cond_1096;
      end 
      if(__stream_matmul_33_stream_ivalid_21 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_104 <= __delay_data_1647__delay_1646__delay_1645___plus_1250;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1860 <= _mul_rshift_round_clip_7_source_start;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1861 <= _tmp_1860;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1862 <= _tmp_1861;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1863 <= _mul_rshift_round_clip_7_source_start;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1864 <= _tmp_1863;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1865 <= _tmp_1864;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1866 <= _tmp_1865;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1867 <= _tmp_1866;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1868 <= _tmp_1867;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1869 <= _tmp_1868;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1870 <= _tmp_1869;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1871 <= _tmp_1870;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1872 <= _tmp_1871;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1873 <= _mul_rshift_round_clip_7_source_stop;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1874 <= _tmp_1873;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1875 <= _tmp_1874;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1876 <= _tmp_1875;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1877 <= _tmp_1876;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1878 <= _tmp_1877;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1879 <= _tmp_1878;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1880 <= _tmp_1879;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1881 <= _tmp_1880;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1882 <= _tmp_1881;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1883 <= _mul_rshift_round_clip_7_source_busy;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1884 <= _tmp_1883;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1885 <= _tmp_1884;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1886 <= _tmp_1885;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1887 <= _tmp_1886;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1888 <= _tmp_1887;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1889 <= _tmp_1888;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1890 <= _tmp_1889;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1891 <= _tmp_1890;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1892 <= _tmp_1891;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1893 <= _mul_rshift_round_clip_7_sink_busy;
      end 
      if(!_mul_rshift_round_clip_7_sink_busy && _tmp_1893) begin
        _mul_rshift_round_clip_7_busy_reg <= 0;
      end 
      if(_mul_rshift_round_clip_7_source_busy) begin
        _mul_rshift_round_clip_7_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_rshift_round_clip_7_fsm_1 = 1;
  localparam _mul_rshift_round_clip_7_fsm_2 = 2;
  localparam _mul_rshift_round_clip_7_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_7_fsm <= _mul_rshift_round_clip_7_fsm_init;
      _mul_rshift_round_clip_7_source_start <= 0;
      _mul_rshift_round_clip_7_source_busy <= 0;
      _mul_rshift_round_clip_7_stream_ivalid <= 0;
    end else begin
      if(__stream_matmul_33_stream_ivalid_21 && _stream_matmul_33_stream_oready) begin
        _mul_rshift_round_clip_7_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_busy) begin
        _mul_rshift_round_clip_7_source_busy <= _stream_matmul_33_source_busy;
      end 
      if(_mul_rshift_round_clip_7_stream_oready && _tmp_1862) begin
        _mul_rshift_round_clip_7_stream_ivalid <= 1;
      end 
      if(_mul_rshift_round_clip_7_stream_oready && 1'd0) begin
        _mul_rshift_round_clip_7_stream_ivalid <= 0;
      end 
      case(_mul_rshift_round_clip_7_fsm)
        _mul_rshift_round_clip_7_fsm_init: begin
          if(_mul_rshift_round_clip_7_run_flag) begin
            _mul_rshift_round_clip_7_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_7_run_flag) begin
            _mul_rshift_round_clip_7_fsm <= _mul_rshift_round_clip_7_fsm_1;
          end 
        end
        _mul_rshift_round_clip_7_fsm_1: begin
          if(_mul_rshift_round_clip_7_source_start && _mul_rshift_round_clip_7_stream_oready) begin
            _mul_rshift_round_clip_7_source_start <= 0;
            _mul_rshift_round_clip_7_source_busy <= 1;
          end 
          if(_mul_rshift_round_clip_7_source_start && _mul_rshift_round_clip_7_stream_oready) begin
            _mul_rshift_round_clip_7_fsm <= _mul_rshift_round_clip_7_fsm_2;
          end 
        end
        _mul_rshift_round_clip_7_fsm_2: begin
          if(_mul_rshift_round_clip_7_stream_oready) begin
            _mul_rshift_round_clip_7_fsm <= _mul_rshift_round_clip_7_fsm_3;
          end 
        end
        _mul_rshift_round_clip_7_fsm_3: begin
          if(_mul_rshift_round_clip_7_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_7_source_busy <= 0;
          end 
          if(_mul_rshift_round_clip_7_stream_oready && 1'd0 && _mul_rshift_round_clip_7_run_flag) begin
            _mul_rshift_round_clip_7_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_7_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_7_fsm <= _mul_rshift_round_clip_7_fsm_init;
          end 
          if(_mul_rshift_round_clip_7_stream_oready && 1'd0 && _mul_rshift_round_clip_7_run_flag) begin
            _mul_rshift_round_clip_7_fsm <= _mul_rshift_round_clip_7_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_8_x_source_ram_renable <= 0;
      _mul_8_x_source_fifo_deq <= 0;
      _mul_8_x_idle <= 1;
      _mul_8_y_source_ram_renable <= 0;
      _mul_8_y_source_fifo_deq <= 0;
      _mul_8_y_idle <= 1;
      _mul_8_rshift_source_ram_renable <= 0;
      _mul_8_rshift_source_fifo_deq <= 0;
      _mul_8_rshift_idle <= 1;
      _mul_8_z_sink_wenable <= 0;
      _mul_8_z_sink_fifo_enq <= 0;
      __mul_8_stream_ivalid_1 <= 0;
      __mul_8_stream_ivalid_2 <= 0;
      __mul_8_stream_ivalid_3 <= 0;
      __mul_8_stream_ivalid_4 <= 0;
      __mul_8_stream_ivalid_5 <= 0;
      __mul_8_stream_ivalid_6 <= 0;
      __mul_8_stream_ivalid_7 <= 0;
      __mul_8_stream_ivalid_8 <= 0;
      _greaterthan_data_139 <= 0;
      _minus_data_141 <= 0;
      _greatereq_data_152 <= 0;
      __delay_data_721__variable_136 <= 0;
      __delay_data_724__variable_137 <= 0;
      __delay_data_727__variable_138 <= 0;
      _sll_data_143 <= 0;
      __delay_data_718_greaterthan_139 <= 0;
      __delay_data_719_greatereq_152 <= 0;
      __delay_data_722__delay_721__variable_136 <= 0;
      __delay_data_725__delay_724__variable_137 <= 0;
      __delay_data_728__delay_727__variable_138 <= 0;
      _cond_data_149 <= 0;
      __delay_data_720__delay_719_greatereq_152 <= 0;
      __delay_data_723__delay_722__delay_721__variable_136 <= 0;
      __delay_data_726__delay_725__delay_724__variable_137 <= 0;
      __delay_data_729__delay_728__delay_727__variable_138 <= 0;
      __muladd_madd_odata_reg_155 <= 0;
      __delay_data_730__delay_729__delay_728____variable_138 <= 0;
      __delay_data_731__delay_730__delay_729____variable_138 <= 0;
      __delay_data_732__delay_731__delay_730____variable_138 <= 0;
      __delay_data_733__delay_732__delay_731____variable_138 <= 0;
      _sra_data_156 <= 0;
      __variable_wdata_136 <= 0;
      __variable_wdata_137 <= 0;
      __variable_wdata_138 <= 0;
      _tmp_629 <= 0;
      _tmp_630 <= 0;
      _tmp_631 <= 0;
      _tmp_632 <= 0;
      _tmp_633 <= 0;
      _tmp_634 <= 0;
      _tmp_635 <= 0;
      _tmp_636 <= 0;
      _tmp_637 <= 0;
      _tmp_638 <= 0;
      _tmp_639 <= 0;
      _tmp_640 <= 0;
      _tmp_641 <= 0;
      _tmp_642 <= 0;
      _tmp_643 <= 0;
      _tmp_644 <= 0;
      _tmp_645 <= 0;
      _tmp_646 <= 0;
      _tmp_647 <= 0;
      _tmp_648 <= 0;
      _tmp_649 <= 0;
      _tmp_650 <= 0;
      _tmp_651 <= 0;
      _tmp_652 <= 0;
      _tmp_653 <= 0;
      _tmp_654 <= 0;
      _tmp_655 <= 0;
      _tmp_656 <= 0;
      _tmp_657 <= 0;
      _tmp_658 <= 0;
      _tmp_659 <= 0;
      _tmp_660 <= 0;
      _tmp_661 <= 0;
      _tmp_662 <= 0;
      _mul_8_busy_reg <= 0;
    end else begin
      if(_mul_8_stream_oready) begin
        _mul_8_x_source_ram_renable <= 0;
        _mul_8_x_source_fifo_deq <= 0;
      end 
      _mul_8_x_idle <= _mul_8_x_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_y_source_ram_renable <= 0;
        _mul_8_y_source_fifo_deq <= 0;
      end 
      _mul_8_y_idle <= _mul_8_y_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_rshift_source_ram_renable <= 0;
        _mul_8_rshift_source_fifo_deq <= 0;
      end 
      _mul_8_rshift_idle <= _mul_8_rshift_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_z_sink_wenable <= 0;
        _mul_8_z_sink_fifo_enq <= 0;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_1 <= _mul_8_stream_ivalid;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_2 <= __mul_8_stream_ivalid_1;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_3 <= __mul_8_stream_ivalid_2;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_4 <= __mul_8_stream_ivalid_3;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_5 <= __mul_8_stream_ivalid_4;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_6 <= __mul_8_stream_ivalid_5;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_7 <= __mul_8_stream_ivalid_6;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_8 <= __mul_8_stream_ivalid_7;
      end 
      if(_mul_8_stream_oready) begin
        _greaterthan_data_139 <= mul_8_rshift_data > 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        _minus_data_141 <= mul_8_rshift_data - 2'sd1;
      end 
      if(_mul_8_stream_oready) begin
        _greatereq_data_152 <= mul_8_x_data >= 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_721__variable_136 <= mul_8_x_data;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_724__variable_137 <= mul_8_y_data;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_727__variable_138 <= mul_8_rshift_data;
      end 
      if(_mul_8_stream_oready) begin
        _sll_data_143 <= 2'sd1 << _minus_data_141;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_718_greaterthan_139 <= _greaterthan_data_139;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_719_greatereq_152 <= _greatereq_data_152;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_722__delay_721__variable_136 <= __delay_data_721__variable_136;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_725__delay_724__variable_137 <= __delay_data_724__variable_137;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_728__delay_727__variable_138 <= __delay_data_727__variable_138;
      end 
      if(_mul_8_stream_oready) begin
        _cond_data_149 <= (__delay_data_718_greaterthan_139)? _sll_data_143 : 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_720__delay_719_greatereq_152 <= __delay_data_719_greatereq_152;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_723__delay_722__delay_721__variable_136 <= __delay_data_722__delay_721__variable_136;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_726__delay_725__delay_724__variable_137 <= __delay_data_725__delay_724__variable_137;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_729__delay_728__delay_727__variable_138 <= __delay_data_728__delay_727__variable_138;
      end 
      if(_mul_8_stream_oready) begin
        __muladd_madd_odata_reg_155 <= __muladd_madd_odata_155;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_730__delay_729__delay_728____variable_138 <= __delay_data_729__delay_728__delay_727__variable_138;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_731__delay_730__delay_729____variable_138 <= __delay_data_730__delay_729__delay_728____variable_138;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_732__delay_731__delay_730____variable_138 <= __delay_data_731__delay_730__delay_729____variable_138;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_733__delay_732__delay_731____variable_138 <= __delay_data_732__delay_731__delay_730____variable_138;
      end 
      if(_mul_8_stream_oready) begin
        _sra_data_156 <= __muladd_data_155 >>> __delay_data_733__delay_732__delay_731____variable_138;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_136 <= _cond_data_700;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_137 <= __delay_data_1264_reinterpretcast_672;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_138 <= _plus_data_734;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_629 <= _mul_8_source_start;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_630 <= _tmp_629;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_631 <= _tmp_630;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_632 <= _mul_8_source_start;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_633 <= _tmp_632;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_634 <= _tmp_633;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_635 <= _tmp_634;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_636 <= _tmp_635;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_637 <= _tmp_636;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_638 <= _tmp_637;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_639 <= _tmp_638;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_640 <= _tmp_639;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_641 <= _tmp_640;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_642 <= _mul_8_source_stop;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_643 <= _tmp_642;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_644 <= _tmp_643;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_645 <= _tmp_644;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_646 <= _tmp_645;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_647 <= _tmp_646;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_648 <= _tmp_647;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_649 <= _tmp_648;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_650 <= _tmp_649;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_651 <= _tmp_650;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_652 <= _mul_8_source_busy;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_653 <= _tmp_652;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_654 <= _tmp_653;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_655 <= _tmp_654;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_656 <= _tmp_655;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_657 <= _tmp_656;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_658 <= _tmp_657;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_659 <= _tmp_658;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_660 <= _tmp_659;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_661 <= _tmp_660;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_662 <= _mul_8_sink_busy;
      end 
      if(!_mul_8_sink_busy && _tmp_662) begin
        _mul_8_busy_reg <= 0;
      end 
      if(_mul_8_source_busy) begin
        _mul_8_busy_reg <= 1;
      end 
      if(__stream_matmul_23_stream_ivalid_1 && _stream_matmul_23_stream_oready) begin
        __variable_wdata_136 <= _cond_data_1033;
      end 
      if(__stream_matmul_23_stream_ivalid_1 && _stream_matmul_23_stream_oready) begin
        __variable_wdata_137 <= __delay_data_1403_reinterpretcast_1029;
      end 
      if(__stream_matmul_23_stream_ivalid_1 && _stream_matmul_23_stream_oready) begin
        __variable_wdata_138 <= _plus_data_1035;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_136 <= _cond_data_1187;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_137 <= _cond_data_1169;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_138 <= __delay_data_1513__delay_1512_plus_1189;
      end 
    end
  end

  localparam _mul_8_fsm_1 = 1;
  localparam _mul_8_fsm_2 = 2;
  localparam _mul_8_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_8_fsm <= _mul_8_fsm_init;
      _mul_8_source_start <= 0;
      _mul_8_source_busy <= 0;
      _mul_8_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_8_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_8_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_8_stream_oready && _tmp_631) begin
        _mul_8_stream_ivalid <= 1;
      end 
      if(_mul_8_stream_oready && 1'd0) begin
        _mul_8_stream_ivalid <= 0;
      end 
      if(__stream_matmul_23_stream_ivalid_1 && _stream_matmul_23_stream_oready) begin
        _mul_8_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_23_stream_oready && _stream_matmul_23_busy) begin
        _mul_8_source_busy <= _stream_matmul_23_source_busy;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        _mul_8_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_busy) begin
        _mul_8_source_busy <= _stream_matmul_33_source_busy;
      end 
      case(_mul_8_fsm)
        _mul_8_fsm_init: begin
          if(_mul_8_run_flag) begin
            _mul_8_source_start <= 1;
          end 
          if(_mul_8_run_flag) begin
            _mul_8_fsm <= _mul_8_fsm_1;
          end 
        end
        _mul_8_fsm_1: begin
          if(_mul_8_source_start && _mul_8_stream_oready) begin
            _mul_8_source_start <= 0;
            _mul_8_source_busy <= 1;
          end 
          if(_mul_8_source_start && _mul_8_stream_oready) begin
            _mul_8_fsm <= _mul_8_fsm_2;
          end 
        end
        _mul_8_fsm_2: begin
          if(_mul_8_stream_oready) begin
            _mul_8_fsm <= _mul_8_fsm_3;
          end 
        end
        _mul_8_fsm_3: begin
          if(_mul_8_stream_oready && 1'd0) begin
            _mul_8_source_busy <= 0;
          end 
          if(_mul_8_stream_oready && 1'd0 && _mul_8_run_flag) begin
            _mul_8_source_start <= 1;
          end 
          if(_mul_8_stream_oready && 1'd0) begin
            _mul_8_fsm <= _mul_8_fsm_init;
          end 
          if(_mul_8_stream_oready && 1'd0 && _mul_8_run_flag) begin
            _mul_8_fsm <= _mul_8_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_9_x_source_ram_renable <= 0;
      _mul_9_x_source_fifo_deq <= 0;
      _mul_9_x_idle <= 1;
      _mul_9_y_source_ram_renable <= 0;
      _mul_9_y_source_fifo_deq <= 0;
      _mul_9_y_idle <= 1;
      _mul_9_rshift_source_ram_renable <= 0;
      _mul_9_rshift_source_fifo_deq <= 0;
      _mul_9_rshift_idle <= 1;
      _mul_9_z_sink_wenable <= 0;
      _mul_9_z_sink_fifo_enq <= 0;
      __mul_9_stream_ivalid_1 <= 0;
      __mul_9_stream_ivalid_2 <= 0;
      __mul_9_stream_ivalid_3 <= 0;
      __mul_9_stream_ivalid_4 <= 0;
      __mul_9_stream_ivalid_5 <= 0;
      __mul_9_stream_ivalid_6 <= 0;
      __mul_9_stream_ivalid_7 <= 0;
      __mul_9_stream_ivalid_8 <= 0;
      _greaterthan_data_160 <= 0;
      _minus_data_162 <= 0;
      _greatereq_data_173 <= 0;
      __delay_data_740__variable_157 <= 0;
      __delay_data_743__variable_158 <= 0;
      __delay_data_746__variable_159 <= 0;
      _sll_data_164 <= 0;
      __delay_data_737_greaterthan_160 <= 0;
      __delay_data_738_greatereq_173 <= 0;
      __delay_data_741__delay_740__variable_157 <= 0;
      __delay_data_744__delay_743__variable_158 <= 0;
      __delay_data_747__delay_746__variable_159 <= 0;
      _cond_data_170 <= 0;
      __delay_data_739__delay_738_greatereq_173 <= 0;
      __delay_data_742__delay_741__delay_740__variable_157 <= 0;
      __delay_data_745__delay_744__delay_743__variable_158 <= 0;
      __delay_data_748__delay_747__delay_746__variable_159 <= 0;
      __muladd_madd_odata_reg_176 <= 0;
      __delay_data_749__delay_748__delay_747____variable_159 <= 0;
      __delay_data_750__delay_749__delay_748____variable_159 <= 0;
      __delay_data_751__delay_750__delay_749____variable_159 <= 0;
      __delay_data_752__delay_751__delay_750____variable_159 <= 0;
      _sra_data_177 <= 0;
      __variable_wdata_157 <= 0;
      __variable_wdata_158 <= 0;
      __variable_wdata_159 <= 0;
      _tmp_663 <= 0;
      _tmp_664 <= 0;
      _tmp_665 <= 0;
      _tmp_666 <= 0;
      _tmp_667 <= 0;
      _tmp_668 <= 0;
      _tmp_669 <= 0;
      _tmp_670 <= 0;
      _tmp_671 <= 0;
      _tmp_672 <= 0;
      _tmp_673 <= 0;
      _tmp_674 <= 0;
      _tmp_675 <= 0;
      _tmp_676 <= 0;
      _tmp_677 <= 0;
      _tmp_678 <= 0;
      _tmp_679 <= 0;
      _tmp_680 <= 0;
      _tmp_681 <= 0;
      _tmp_682 <= 0;
      _tmp_683 <= 0;
      _tmp_684 <= 0;
      _tmp_685 <= 0;
      _tmp_686 <= 0;
      _tmp_687 <= 0;
      _tmp_688 <= 0;
      _tmp_689 <= 0;
      _tmp_690 <= 0;
      _tmp_691 <= 0;
      _tmp_692 <= 0;
      _tmp_693 <= 0;
      _tmp_694 <= 0;
      _tmp_695 <= 0;
      _tmp_696 <= 0;
      _mul_9_busy_reg <= 0;
    end else begin
      if(_mul_9_stream_oready) begin
        _mul_9_x_source_ram_renable <= 0;
        _mul_9_x_source_fifo_deq <= 0;
      end 
      _mul_9_x_idle <= _mul_9_x_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_y_source_ram_renable <= 0;
        _mul_9_y_source_fifo_deq <= 0;
      end 
      _mul_9_y_idle <= _mul_9_y_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_rshift_source_ram_renable <= 0;
        _mul_9_rshift_source_fifo_deq <= 0;
      end 
      _mul_9_rshift_idle <= _mul_9_rshift_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_z_sink_wenable <= 0;
        _mul_9_z_sink_fifo_enq <= 0;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_1 <= _mul_9_stream_ivalid;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_2 <= __mul_9_stream_ivalid_1;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_3 <= __mul_9_stream_ivalid_2;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_4 <= __mul_9_stream_ivalid_3;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_5 <= __mul_9_stream_ivalid_4;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_6 <= __mul_9_stream_ivalid_5;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_7 <= __mul_9_stream_ivalid_6;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_8 <= __mul_9_stream_ivalid_7;
      end 
      if(_mul_9_stream_oready) begin
        _greaterthan_data_160 <= mul_9_rshift_data > 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        _minus_data_162 <= mul_9_rshift_data - 2'sd1;
      end 
      if(_mul_9_stream_oready) begin
        _greatereq_data_173 <= mul_9_x_data >= 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_740__variable_157 <= mul_9_x_data;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_743__variable_158 <= mul_9_y_data;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_746__variable_159 <= mul_9_rshift_data;
      end 
      if(_mul_9_stream_oready) begin
        _sll_data_164 <= 2'sd1 << _minus_data_162;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_737_greaterthan_160 <= _greaterthan_data_160;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_738_greatereq_173 <= _greatereq_data_173;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_741__delay_740__variable_157 <= __delay_data_740__variable_157;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_744__delay_743__variable_158 <= __delay_data_743__variable_158;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_747__delay_746__variable_159 <= __delay_data_746__variable_159;
      end 
      if(_mul_9_stream_oready) begin
        _cond_data_170 <= (__delay_data_737_greaterthan_160)? _sll_data_164 : 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_739__delay_738_greatereq_173 <= __delay_data_738_greatereq_173;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_742__delay_741__delay_740__variable_157 <= __delay_data_741__delay_740__variable_157;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_745__delay_744__delay_743__variable_158 <= __delay_data_744__delay_743__variable_158;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_748__delay_747__delay_746__variable_159 <= __delay_data_747__delay_746__variable_159;
      end 
      if(_mul_9_stream_oready) begin
        __muladd_madd_odata_reg_176 <= __muladd_madd_odata_176;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_749__delay_748__delay_747____variable_159 <= __delay_data_748__delay_747__delay_746__variable_159;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_750__delay_749__delay_748____variable_159 <= __delay_data_749__delay_748__delay_747____variable_159;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_751__delay_750__delay_749____variable_159 <= __delay_data_750__delay_749__delay_748____variable_159;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_752__delay_751__delay_750____variable_159 <= __delay_data_751__delay_750__delay_749____variable_159;
      end 
      if(_mul_9_stream_oready) begin
        _sra_data_177 <= __muladd_data_176 >>> __delay_data_752__delay_751__delay_750____variable_159;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_157 <= _cond_data_702;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_158 <= __delay_data_1266_reinterpretcast_673;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_159 <= _plus_data_753;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_663 <= _mul_9_source_start;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_664 <= _tmp_663;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_665 <= _tmp_664;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_666 <= _mul_9_source_start;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_667 <= _tmp_666;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_668 <= _tmp_667;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_669 <= _tmp_668;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_670 <= _tmp_669;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_671 <= _tmp_670;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_672 <= _tmp_671;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_673 <= _tmp_672;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_674 <= _tmp_673;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_675 <= _tmp_674;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_676 <= _mul_9_source_stop;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_677 <= _tmp_676;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_678 <= _tmp_677;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_679 <= _tmp_678;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_680 <= _tmp_679;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_681 <= _tmp_680;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_682 <= _tmp_681;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_683 <= _tmp_682;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_684 <= _tmp_683;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_685 <= _tmp_684;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_686 <= _mul_9_source_busy;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_687 <= _tmp_686;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_688 <= _tmp_687;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_689 <= _tmp_688;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_690 <= _tmp_689;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_691 <= _tmp_690;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_692 <= _tmp_691;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_693 <= _tmp_692;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_694 <= _tmp_693;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_695 <= _tmp_694;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_696 <= _mul_9_sink_busy;
      end 
      if(!_mul_9_sink_busy && _tmp_696) begin
        _mul_9_busy_reg <= 0;
      end 
      if(_mul_9_source_busy) begin
        _mul_9_busy_reg <= 1;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_157 <= _cond_data_1192;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_158 <= _cond_data_1171;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_159 <= __delay_data_1522__delay_1521_plus_1194;
      end 
    end
  end

  localparam _mul_9_fsm_1 = 1;
  localparam _mul_9_fsm_2 = 2;
  localparam _mul_9_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_9_fsm <= _mul_9_fsm_init;
      _mul_9_source_start <= 0;
      _mul_9_source_busy <= 0;
      _mul_9_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_9_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_9_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_9_stream_oready && _tmp_665) begin
        _mul_9_stream_ivalid <= 1;
      end 
      if(_mul_9_stream_oready && 1'd0) begin
        _mul_9_stream_ivalid <= 0;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        _mul_9_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_busy) begin
        _mul_9_source_busy <= _stream_matmul_33_source_busy;
      end 
      case(_mul_9_fsm)
        _mul_9_fsm_init: begin
          if(_mul_9_run_flag) begin
            _mul_9_source_start <= 1;
          end 
          if(_mul_9_run_flag) begin
            _mul_9_fsm <= _mul_9_fsm_1;
          end 
        end
        _mul_9_fsm_1: begin
          if(_mul_9_source_start && _mul_9_stream_oready) begin
            _mul_9_source_start <= 0;
            _mul_9_source_busy <= 1;
          end 
          if(_mul_9_source_start && _mul_9_stream_oready) begin
            _mul_9_fsm <= _mul_9_fsm_2;
          end 
        end
        _mul_9_fsm_2: begin
          if(_mul_9_stream_oready) begin
            _mul_9_fsm <= _mul_9_fsm_3;
          end 
        end
        _mul_9_fsm_3: begin
          if(_mul_9_stream_oready && 1'd0) begin
            _mul_9_source_busy <= 0;
          end 
          if(_mul_9_stream_oready && 1'd0 && _mul_9_run_flag) begin
            _mul_9_source_start <= 1;
          end 
          if(_mul_9_stream_oready && 1'd0) begin
            _mul_9_fsm <= _mul_9_fsm_init;
          end 
          if(_mul_9_stream_oready && 1'd0 && _mul_9_run_flag) begin
            _mul_9_fsm <= _mul_9_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_10_x_source_ram_renable <= 0;
      _mul_10_x_source_fifo_deq <= 0;
      _mul_10_x_idle <= 1;
      _mul_10_y_source_ram_renable <= 0;
      _mul_10_y_source_fifo_deq <= 0;
      _mul_10_y_idle <= 1;
      _mul_10_rshift_source_ram_renable <= 0;
      _mul_10_rshift_source_fifo_deq <= 0;
      _mul_10_rshift_idle <= 1;
      _mul_10_z_sink_wenable <= 0;
      _mul_10_z_sink_fifo_enq <= 0;
      __mul_10_stream_ivalid_1 <= 0;
      __mul_10_stream_ivalid_2 <= 0;
      __mul_10_stream_ivalid_3 <= 0;
      __mul_10_stream_ivalid_4 <= 0;
      __mul_10_stream_ivalid_5 <= 0;
      __mul_10_stream_ivalid_6 <= 0;
      __mul_10_stream_ivalid_7 <= 0;
      __mul_10_stream_ivalid_8 <= 0;
      _greaterthan_data_181 <= 0;
      _minus_data_183 <= 0;
      _greatereq_data_194 <= 0;
      __delay_data_759__variable_178 <= 0;
      __delay_data_762__variable_179 <= 0;
      __delay_data_765__variable_180 <= 0;
      _sll_data_185 <= 0;
      __delay_data_756_greaterthan_181 <= 0;
      __delay_data_757_greatereq_194 <= 0;
      __delay_data_760__delay_759__variable_178 <= 0;
      __delay_data_763__delay_762__variable_179 <= 0;
      __delay_data_766__delay_765__variable_180 <= 0;
      _cond_data_191 <= 0;
      __delay_data_758__delay_757_greatereq_194 <= 0;
      __delay_data_761__delay_760__delay_759__variable_178 <= 0;
      __delay_data_764__delay_763__delay_762__variable_179 <= 0;
      __delay_data_767__delay_766__delay_765__variable_180 <= 0;
      __muladd_madd_odata_reg_197 <= 0;
      __delay_data_768__delay_767__delay_766____variable_180 <= 0;
      __delay_data_769__delay_768__delay_767____variable_180 <= 0;
      __delay_data_770__delay_769__delay_768____variable_180 <= 0;
      __delay_data_771__delay_770__delay_769____variable_180 <= 0;
      _sra_data_198 <= 0;
      __variable_wdata_178 <= 0;
      __variable_wdata_179 <= 0;
      __variable_wdata_180 <= 0;
      _tmp_697 <= 0;
      _tmp_698 <= 0;
      _tmp_699 <= 0;
      _tmp_700 <= 0;
      _tmp_701 <= 0;
      _tmp_702 <= 0;
      _tmp_703 <= 0;
      _tmp_704 <= 0;
      _tmp_705 <= 0;
      _tmp_706 <= 0;
      _tmp_707 <= 0;
      _tmp_708 <= 0;
      _tmp_709 <= 0;
      _tmp_710 <= 0;
      _tmp_711 <= 0;
      _tmp_712 <= 0;
      _tmp_713 <= 0;
      _tmp_714 <= 0;
      _tmp_715 <= 0;
      _tmp_716 <= 0;
      _tmp_717 <= 0;
      _tmp_718 <= 0;
      _tmp_719 <= 0;
      _tmp_720 <= 0;
      _tmp_721 <= 0;
      _tmp_722 <= 0;
      _tmp_723 <= 0;
      _tmp_724 <= 0;
      _tmp_725 <= 0;
      _tmp_726 <= 0;
      _tmp_727 <= 0;
      _tmp_728 <= 0;
      _tmp_729 <= 0;
      _tmp_730 <= 0;
      _mul_10_busy_reg <= 0;
    end else begin
      if(_mul_10_stream_oready) begin
        _mul_10_x_source_ram_renable <= 0;
        _mul_10_x_source_fifo_deq <= 0;
      end 
      _mul_10_x_idle <= _mul_10_x_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_y_source_ram_renable <= 0;
        _mul_10_y_source_fifo_deq <= 0;
      end 
      _mul_10_y_idle <= _mul_10_y_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_rshift_source_ram_renable <= 0;
        _mul_10_rshift_source_fifo_deq <= 0;
      end 
      _mul_10_rshift_idle <= _mul_10_rshift_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_z_sink_wenable <= 0;
        _mul_10_z_sink_fifo_enq <= 0;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_1 <= _mul_10_stream_ivalid;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_2 <= __mul_10_stream_ivalid_1;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_3 <= __mul_10_stream_ivalid_2;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_4 <= __mul_10_stream_ivalid_3;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_5 <= __mul_10_stream_ivalid_4;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_6 <= __mul_10_stream_ivalid_5;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_7 <= __mul_10_stream_ivalid_6;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_8 <= __mul_10_stream_ivalid_7;
      end 
      if(_mul_10_stream_oready) begin
        _greaterthan_data_181 <= mul_10_rshift_data > 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        _minus_data_183 <= mul_10_rshift_data - 2'sd1;
      end 
      if(_mul_10_stream_oready) begin
        _greatereq_data_194 <= mul_10_x_data >= 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_759__variable_178 <= mul_10_x_data;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_762__variable_179 <= mul_10_y_data;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_765__variable_180 <= mul_10_rshift_data;
      end 
      if(_mul_10_stream_oready) begin
        _sll_data_185 <= 2'sd1 << _minus_data_183;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_756_greaterthan_181 <= _greaterthan_data_181;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_757_greatereq_194 <= _greatereq_data_194;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_760__delay_759__variable_178 <= __delay_data_759__variable_178;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_763__delay_762__variable_179 <= __delay_data_762__variable_179;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_766__delay_765__variable_180 <= __delay_data_765__variable_180;
      end 
      if(_mul_10_stream_oready) begin
        _cond_data_191 <= (__delay_data_756_greaterthan_181)? _sll_data_185 : 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_758__delay_757_greatereq_194 <= __delay_data_757_greatereq_194;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_761__delay_760__delay_759__variable_178 <= __delay_data_760__delay_759__variable_178;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_764__delay_763__delay_762__variable_179 <= __delay_data_763__delay_762__variable_179;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_767__delay_766__delay_765__variable_180 <= __delay_data_766__delay_765__variable_180;
      end 
      if(_mul_10_stream_oready) begin
        __muladd_madd_odata_reg_197 <= __muladd_madd_odata_197;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_768__delay_767__delay_766____variable_180 <= __delay_data_767__delay_766__delay_765__variable_180;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_769__delay_768__delay_767____variable_180 <= __delay_data_768__delay_767__delay_766____variable_180;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_770__delay_769__delay_768____variable_180 <= __delay_data_769__delay_768__delay_767____variable_180;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_771__delay_770__delay_769____variable_180 <= __delay_data_770__delay_769__delay_768____variable_180;
      end 
      if(_mul_10_stream_oready) begin
        _sra_data_198 <= __muladd_data_197 >>> __delay_data_771__delay_770__delay_769____variable_180;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_178 <= _cond_data_704;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_179 <= __delay_data_1268_reinterpretcast_674;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_180 <= _plus_data_772;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_697 <= _mul_10_source_start;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_698 <= _tmp_697;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_699 <= _tmp_698;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_700 <= _mul_10_source_start;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_701 <= _tmp_700;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_702 <= _tmp_701;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_703 <= _tmp_702;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_704 <= _tmp_703;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_705 <= _tmp_704;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_706 <= _tmp_705;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_707 <= _tmp_706;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_708 <= _tmp_707;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_709 <= _tmp_708;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_710 <= _mul_10_source_stop;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_711 <= _tmp_710;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_712 <= _tmp_711;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_713 <= _tmp_712;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_714 <= _tmp_713;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_715 <= _tmp_714;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_716 <= _tmp_715;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_717 <= _tmp_716;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_718 <= _tmp_717;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_719 <= _tmp_718;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_720 <= _mul_10_source_busy;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_721 <= _tmp_720;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_722 <= _tmp_721;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_723 <= _tmp_722;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_724 <= _tmp_723;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_725 <= _tmp_724;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_726 <= _tmp_725;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_727 <= _tmp_726;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_728 <= _tmp_727;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_729 <= _tmp_728;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_730 <= _mul_10_sink_busy;
      end 
      if(!_mul_10_sink_busy && _tmp_730) begin
        _mul_10_busy_reg <= 0;
      end 
      if(_mul_10_source_busy) begin
        _mul_10_busy_reg <= 1;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_178 <= _cond_data_1208;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_179 <= _cond_data_1181;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_180 <= __delay_data_1568__delay_1567_plus_1210;
      end 
    end
  end

  localparam _mul_10_fsm_1 = 1;
  localparam _mul_10_fsm_2 = 2;
  localparam _mul_10_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_10_fsm <= _mul_10_fsm_init;
      _mul_10_source_start <= 0;
      _mul_10_source_busy <= 0;
      _mul_10_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_10_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_10_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_10_stream_oready && _tmp_699) begin
        _mul_10_stream_ivalid <= 1;
      end 
      if(_mul_10_stream_oready && 1'd0) begin
        _mul_10_stream_ivalid <= 0;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        _mul_10_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_busy) begin
        _mul_10_source_busy <= _stream_matmul_33_source_busy;
      end 
      case(_mul_10_fsm)
        _mul_10_fsm_init: begin
          if(_mul_10_run_flag) begin
            _mul_10_source_start <= 1;
          end 
          if(_mul_10_run_flag) begin
            _mul_10_fsm <= _mul_10_fsm_1;
          end 
        end
        _mul_10_fsm_1: begin
          if(_mul_10_source_start && _mul_10_stream_oready) begin
            _mul_10_source_start <= 0;
            _mul_10_source_busy <= 1;
          end 
          if(_mul_10_source_start && _mul_10_stream_oready) begin
            _mul_10_fsm <= _mul_10_fsm_2;
          end 
        end
        _mul_10_fsm_2: begin
          if(_mul_10_stream_oready) begin
            _mul_10_fsm <= _mul_10_fsm_3;
          end 
        end
        _mul_10_fsm_3: begin
          if(_mul_10_stream_oready && 1'd0) begin
            _mul_10_source_busy <= 0;
          end 
          if(_mul_10_stream_oready && 1'd0 && _mul_10_run_flag) begin
            _mul_10_source_start <= 1;
          end 
          if(_mul_10_stream_oready && 1'd0) begin
            _mul_10_fsm <= _mul_10_fsm_init;
          end 
          if(_mul_10_stream_oready && 1'd0 && _mul_10_run_flag) begin
            _mul_10_fsm <= _mul_10_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_11_x_source_ram_renable <= 0;
      _mul_11_x_source_fifo_deq <= 0;
      _mul_11_x_idle <= 1;
      _mul_11_y_source_ram_renable <= 0;
      _mul_11_y_source_fifo_deq <= 0;
      _mul_11_y_idle <= 1;
      _mul_11_rshift_source_ram_renable <= 0;
      _mul_11_rshift_source_fifo_deq <= 0;
      _mul_11_rshift_idle <= 1;
      _mul_11_z_sink_wenable <= 0;
      _mul_11_z_sink_fifo_enq <= 0;
      __mul_11_stream_ivalid_1 <= 0;
      __mul_11_stream_ivalid_2 <= 0;
      __mul_11_stream_ivalid_3 <= 0;
      __mul_11_stream_ivalid_4 <= 0;
      __mul_11_stream_ivalid_5 <= 0;
      __mul_11_stream_ivalid_6 <= 0;
      __mul_11_stream_ivalid_7 <= 0;
      __mul_11_stream_ivalid_8 <= 0;
      _greaterthan_data_202 <= 0;
      _minus_data_204 <= 0;
      _greatereq_data_215 <= 0;
      __delay_data_778__variable_199 <= 0;
      __delay_data_781__variable_200 <= 0;
      __delay_data_784__variable_201 <= 0;
      _sll_data_206 <= 0;
      __delay_data_775_greaterthan_202 <= 0;
      __delay_data_776_greatereq_215 <= 0;
      __delay_data_779__delay_778__variable_199 <= 0;
      __delay_data_782__delay_781__variable_200 <= 0;
      __delay_data_785__delay_784__variable_201 <= 0;
      _cond_data_212 <= 0;
      __delay_data_777__delay_776_greatereq_215 <= 0;
      __delay_data_780__delay_779__delay_778__variable_199 <= 0;
      __delay_data_783__delay_782__delay_781__variable_200 <= 0;
      __delay_data_786__delay_785__delay_784__variable_201 <= 0;
      __muladd_madd_odata_reg_218 <= 0;
      __delay_data_787__delay_786__delay_785____variable_201 <= 0;
      __delay_data_788__delay_787__delay_786____variable_201 <= 0;
      __delay_data_789__delay_788__delay_787____variable_201 <= 0;
      __delay_data_790__delay_789__delay_788____variable_201 <= 0;
      _sra_data_219 <= 0;
      __variable_wdata_199 <= 0;
      __variable_wdata_200 <= 0;
      __variable_wdata_201 <= 0;
      _tmp_731 <= 0;
      _tmp_732 <= 0;
      _tmp_733 <= 0;
      _tmp_734 <= 0;
      _tmp_735 <= 0;
      _tmp_736 <= 0;
      _tmp_737 <= 0;
      _tmp_738 <= 0;
      _tmp_739 <= 0;
      _tmp_740 <= 0;
      _tmp_741 <= 0;
      _tmp_742 <= 0;
      _tmp_743 <= 0;
      _tmp_744 <= 0;
      _tmp_745 <= 0;
      _tmp_746 <= 0;
      _tmp_747 <= 0;
      _tmp_748 <= 0;
      _tmp_749 <= 0;
      _tmp_750 <= 0;
      _tmp_751 <= 0;
      _tmp_752 <= 0;
      _tmp_753 <= 0;
      _tmp_754 <= 0;
      _tmp_755 <= 0;
      _tmp_756 <= 0;
      _tmp_757 <= 0;
      _tmp_758 <= 0;
      _tmp_759 <= 0;
      _tmp_760 <= 0;
      _tmp_761 <= 0;
      _tmp_762 <= 0;
      _tmp_763 <= 0;
      _tmp_764 <= 0;
      _mul_11_busy_reg <= 0;
    end else begin
      if(_mul_11_stream_oready) begin
        _mul_11_x_source_ram_renable <= 0;
        _mul_11_x_source_fifo_deq <= 0;
      end 
      _mul_11_x_idle <= _mul_11_x_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_y_source_ram_renable <= 0;
        _mul_11_y_source_fifo_deq <= 0;
      end 
      _mul_11_y_idle <= _mul_11_y_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_rshift_source_ram_renable <= 0;
        _mul_11_rshift_source_fifo_deq <= 0;
      end 
      _mul_11_rshift_idle <= _mul_11_rshift_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_z_sink_wenable <= 0;
        _mul_11_z_sink_fifo_enq <= 0;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_1 <= _mul_11_stream_ivalid;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_2 <= __mul_11_stream_ivalid_1;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_3 <= __mul_11_stream_ivalid_2;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_4 <= __mul_11_stream_ivalid_3;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_5 <= __mul_11_stream_ivalid_4;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_6 <= __mul_11_stream_ivalid_5;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_7 <= __mul_11_stream_ivalid_6;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_8 <= __mul_11_stream_ivalid_7;
      end 
      if(_mul_11_stream_oready) begin
        _greaterthan_data_202 <= mul_11_rshift_data > 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        _minus_data_204 <= mul_11_rshift_data - 2'sd1;
      end 
      if(_mul_11_stream_oready) begin
        _greatereq_data_215 <= mul_11_x_data >= 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_778__variable_199 <= mul_11_x_data;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_781__variable_200 <= mul_11_y_data;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_784__variable_201 <= mul_11_rshift_data;
      end 
      if(_mul_11_stream_oready) begin
        _sll_data_206 <= 2'sd1 << _minus_data_204;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_775_greaterthan_202 <= _greaterthan_data_202;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_776_greatereq_215 <= _greatereq_data_215;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_779__delay_778__variable_199 <= __delay_data_778__variable_199;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_782__delay_781__variable_200 <= __delay_data_781__variable_200;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_785__delay_784__variable_201 <= __delay_data_784__variable_201;
      end 
      if(_mul_11_stream_oready) begin
        _cond_data_212 <= (__delay_data_775_greaterthan_202)? _sll_data_206 : 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_777__delay_776_greatereq_215 <= __delay_data_776_greatereq_215;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_780__delay_779__delay_778__variable_199 <= __delay_data_779__delay_778__variable_199;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_783__delay_782__delay_781__variable_200 <= __delay_data_782__delay_781__variable_200;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_786__delay_785__delay_784__variable_201 <= __delay_data_785__delay_784__variable_201;
      end 
      if(_mul_11_stream_oready) begin
        __muladd_madd_odata_reg_218 <= __muladd_madd_odata_218;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_787__delay_786__delay_785____variable_201 <= __delay_data_786__delay_785__delay_784__variable_201;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_788__delay_787__delay_786____variable_201 <= __delay_data_787__delay_786__delay_785____variable_201;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_789__delay_788__delay_787____variable_201 <= __delay_data_788__delay_787__delay_786____variable_201;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_790__delay_789__delay_788____variable_201 <= __delay_data_789__delay_788__delay_787____variable_201;
      end 
      if(_mul_11_stream_oready) begin
        _sra_data_219 <= __muladd_data_218 >>> __delay_data_790__delay_789__delay_788____variable_201;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_199 <= _cond_data_706;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_200 <= __delay_data_1270_reinterpretcast_675;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_201 <= _plus_data_791;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_731 <= _mul_11_source_start;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_732 <= _tmp_731;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_733 <= _tmp_732;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_734 <= _mul_11_source_start;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_735 <= _tmp_734;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_736 <= _tmp_735;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_737 <= _tmp_736;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_738 <= _tmp_737;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_739 <= _tmp_738;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_740 <= _tmp_739;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_741 <= _tmp_740;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_742 <= _tmp_741;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_743 <= _tmp_742;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_744 <= _mul_11_source_stop;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_745 <= _tmp_744;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_746 <= _tmp_745;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_747 <= _tmp_746;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_748 <= _tmp_747;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_749 <= _tmp_748;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_750 <= _tmp_749;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_751 <= _tmp_750;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_752 <= _tmp_751;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_753 <= _tmp_752;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_754 <= _mul_11_source_busy;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_755 <= _tmp_754;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_756 <= _tmp_755;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_757 <= _tmp_756;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_758 <= _tmp_757;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_759 <= _tmp_758;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_760 <= _tmp_759;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_761 <= _tmp_760;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_762 <= _tmp_761;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_763 <= _tmp_762;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_764 <= _mul_11_sink_busy;
      end 
      if(!_mul_11_sink_busy && _tmp_764) begin
        _mul_11_busy_reg <= 0;
      end 
      if(_mul_11_source_busy) begin
        _mul_11_busy_reg <= 1;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_199 <= _cond_data_1213;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_200 <= _cond_data_1183;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        __variable_wdata_201 <= __delay_data_1573__delay_1572_plus_1215;
      end 
    end
  end

  localparam _mul_11_fsm_1 = 1;
  localparam _mul_11_fsm_2 = 2;
  localparam _mul_11_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_11_fsm <= _mul_11_fsm_init;
      _mul_11_source_start <= 0;
      _mul_11_source_busy <= 0;
      _mul_11_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_11_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_11_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_11_stream_oready && _tmp_733) begin
        _mul_11_stream_ivalid <= 1;
      end 
      if(_mul_11_stream_oready && 1'd0) begin
        _mul_11_stream_ivalid <= 0;
      end 
      if(__stream_matmul_33_stream_ivalid_3 && _stream_matmul_33_stream_oready) begin
        _mul_11_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_busy) begin
        _mul_11_source_busy <= _stream_matmul_33_source_busy;
      end 
      case(_mul_11_fsm)
        _mul_11_fsm_init: begin
          if(_mul_11_run_flag) begin
            _mul_11_source_start <= 1;
          end 
          if(_mul_11_run_flag) begin
            _mul_11_fsm <= _mul_11_fsm_1;
          end 
        end
        _mul_11_fsm_1: begin
          if(_mul_11_source_start && _mul_11_stream_oready) begin
            _mul_11_source_start <= 0;
            _mul_11_source_busy <= 1;
          end 
          if(_mul_11_source_start && _mul_11_stream_oready) begin
            _mul_11_fsm <= _mul_11_fsm_2;
          end 
        end
        _mul_11_fsm_2: begin
          if(_mul_11_stream_oready) begin
            _mul_11_fsm <= _mul_11_fsm_3;
          end 
        end
        _mul_11_fsm_3: begin
          if(_mul_11_stream_oready && 1'd0) begin
            _mul_11_source_busy <= 0;
          end 
          if(_mul_11_stream_oready && 1'd0 && _mul_11_run_flag) begin
            _mul_11_source_start <= 1;
          end 
          if(_mul_11_stream_oready && 1'd0) begin
            _mul_11_fsm <= _mul_11_fsm_init;
          end 
          if(_mul_11_stream_oready && 1'd0 && _mul_11_run_flag) begin
            _mul_11_fsm <= _mul_11_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_12_x_source_ram_renable <= 0;
      _mul_12_x_source_fifo_deq <= 0;
      _mul_12_x_idle <= 1;
      _mul_12_y_source_ram_renable <= 0;
      _mul_12_y_source_fifo_deq <= 0;
      _mul_12_y_idle <= 1;
      _mul_12_rshift_source_ram_renable <= 0;
      _mul_12_rshift_source_fifo_deq <= 0;
      _mul_12_rshift_idle <= 1;
      _mul_12_z_sink_wenable <= 0;
      _mul_12_z_sink_fifo_enq <= 0;
      __mul_12_stream_ivalid_1 <= 0;
      __mul_12_stream_ivalid_2 <= 0;
      __mul_12_stream_ivalid_3 <= 0;
      __mul_12_stream_ivalid_4 <= 0;
      __mul_12_stream_ivalid_5 <= 0;
      __mul_12_stream_ivalid_6 <= 0;
      __mul_12_stream_ivalid_7 <= 0;
      __mul_12_stream_ivalid_8 <= 0;
      _greaterthan_data_223 <= 0;
      _minus_data_225 <= 0;
      _greatereq_data_236 <= 0;
      __delay_data_797__variable_220 <= 0;
      __delay_data_800__variable_221 <= 0;
      __delay_data_803__variable_222 <= 0;
      _sll_data_227 <= 0;
      __delay_data_794_greaterthan_223 <= 0;
      __delay_data_795_greatereq_236 <= 0;
      __delay_data_798__delay_797__variable_220 <= 0;
      __delay_data_801__delay_800__variable_221 <= 0;
      __delay_data_804__delay_803__variable_222 <= 0;
      _cond_data_233 <= 0;
      __delay_data_796__delay_795_greatereq_236 <= 0;
      __delay_data_799__delay_798__delay_797__variable_220 <= 0;
      __delay_data_802__delay_801__delay_800__variable_221 <= 0;
      __delay_data_805__delay_804__delay_803__variable_222 <= 0;
      __muladd_madd_odata_reg_239 <= 0;
      __delay_data_806__delay_805__delay_804____variable_222 <= 0;
      __delay_data_807__delay_806__delay_805____variable_222 <= 0;
      __delay_data_808__delay_807__delay_806____variable_222 <= 0;
      __delay_data_809__delay_808__delay_807____variable_222 <= 0;
      _sra_data_240 <= 0;
      __variable_wdata_220 <= 0;
      __variable_wdata_221 <= 0;
      __variable_wdata_222 <= 0;
      _tmp_765 <= 0;
      _tmp_766 <= 0;
      _tmp_767 <= 0;
      _tmp_768 <= 0;
      _tmp_769 <= 0;
      _tmp_770 <= 0;
      _tmp_771 <= 0;
      _tmp_772 <= 0;
      _tmp_773 <= 0;
      _tmp_774 <= 0;
      _tmp_775 <= 0;
      _tmp_776 <= 0;
      _tmp_777 <= 0;
      _tmp_778 <= 0;
      _tmp_779 <= 0;
      _tmp_780 <= 0;
      _tmp_781 <= 0;
      _tmp_782 <= 0;
      _tmp_783 <= 0;
      _tmp_784 <= 0;
      _tmp_785 <= 0;
      _tmp_786 <= 0;
      _tmp_787 <= 0;
      _tmp_788 <= 0;
      _tmp_789 <= 0;
      _tmp_790 <= 0;
      _tmp_791 <= 0;
      _tmp_792 <= 0;
      _tmp_793 <= 0;
      _tmp_794 <= 0;
      _tmp_795 <= 0;
      _tmp_796 <= 0;
      _tmp_797 <= 0;
      _tmp_798 <= 0;
      _mul_12_busy_reg <= 0;
    end else begin
      if(_mul_12_stream_oready) begin
        _mul_12_x_source_ram_renable <= 0;
        _mul_12_x_source_fifo_deq <= 0;
      end 
      _mul_12_x_idle <= _mul_12_x_idle;
      if(_mul_12_stream_oready) begin
        _mul_12_y_source_ram_renable <= 0;
        _mul_12_y_source_fifo_deq <= 0;
      end 
      _mul_12_y_idle <= _mul_12_y_idle;
      if(_mul_12_stream_oready) begin
        _mul_12_rshift_source_ram_renable <= 0;
        _mul_12_rshift_source_fifo_deq <= 0;
      end 
      _mul_12_rshift_idle <= _mul_12_rshift_idle;
      if(_mul_12_stream_oready) begin
        _mul_12_z_sink_wenable <= 0;
        _mul_12_z_sink_fifo_enq <= 0;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_1 <= _mul_12_stream_ivalid;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_2 <= __mul_12_stream_ivalid_1;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_3 <= __mul_12_stream_ivalid_2;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_4 <= __mul_12_stream_ivalid_3;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_5 <= __mul_12_stream_ivalid_4;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_6 <= __mul_12_stream_ivalid_5;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_7 <= __mul_12_stream_ivalid_6;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_8 <= __mul_12_stream_ivalid_7;
      end 
      if(_mul_12_stream_oready) begin
        _greaterthan_data_223 <= mul_12_rshift_data > 1'sd0;
      end 
      if(_mul_12_stream_oready) begin
        _minus_data_225 <= mul_12_rshift_data - 2'sd1;
      end 
      if(_mul_12_stream_oready) begin
        _greatereq_data_236 <= mul_12_x_data >= 1'sd0;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_797__variable_220 <= mul_12_x_data;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_800__variable_221 <= mul_12_y_data;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_803__variable_222 <= mul_12_rshift_data;
      end 
      if(_mul_12_stream_oready) begin
        _sll_data_227 <= 2'sd1 << _minus_data_225;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_794_greaterthan_223 <= _greaterthan_data_223;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_795_greatereq_236 <= _greatereq_data_236;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_798__delay_797__variable_220 <= __delay_data_797__variable_220;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_801__delay_800__variable_221 <= __delay_data_800__variable_221;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_804__delay_803__variable_222 <= __delay_data_803__variable_222;
      end 
      if(_mul_12_stream_oready) begin
        _cond_data_233 <= (__delay_data_794_greaterthan_223)? _sll_data_227 : 1'sd0;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_796__delay_795_greatereq_236 <= __delay_data_795_greatereq_236;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_799__delay_798__delay_797__variable_220 <= __delay_data_798__delay_797__variable_220;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_802__delay_801__delay_800__variable_221 <= __delay_data_801__delay_800__variable_221;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_805__delay_804__delay_803__variable_222 <= __delay_data_804__delay_803__variable_222;
      end 
      if(_mul_12_stream_oready) begin
        __muladd_madd_odata_reg_239 <= __muladd_madd_odata_239;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_806__delay_805__delay_804____variable_222 <= __delay_data_805__delay_804__delay_803__variable_222;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_807__delay_806__delay_805____variable_222 <= __delay_data_806__delay_805__delay_804____variable_222;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_808__delay_807__delay_806____variable_222 <= __delay_data_807__delay_806__delay_805____variable_222;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_809__delay_808__delay_807____variable_222 <= __delay_data_808__delay_807__delay_806____variable_222;
      end 
      if(_mul_12_stream_oready) begin
        _sra_data_240 <= __muladd_data_239 >>> __delay_data_809__delay_808__delay_807____variable_222;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_220 <= _cond_data_708;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_221 <= __delay_data_1272_reinterpretcast_676;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_222 <= _plus_data_810;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_765 <= _mul_12_source_start;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_766 <= _tmp_765;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_767 <= _tmp_766;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_768 <= _mul_12_source_start;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_769 <= _tmp_768;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_770 <= _tmp_769;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_771 <= _tmp_770;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_772 <= _tmp_771;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_773 <= _tmp_772;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_774 <= _tmp_773;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_775 <= _tmp_774;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_776 <= _tmp_775;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_777 <= _tmp_776;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_778 <= _mul_12_source_stop;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_779 <= _tmp_778;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_780 <= _tmp_779;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_781 <= _tmp_780;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_782 <= _tmp_781;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_783 <= _tmp_782;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_784 <= _tmp_783;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_785 <= _tmp_784;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_786 <= _tmp_785;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_787 <= _tmp_786;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_788 <= _mul_12_source_busy;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_789 <= _tmp_788;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_790 <= _tmp_789;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_791 <= _tmp_790;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_792 <= _tmp_791;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_793 <= _tmp_792;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_794 <= _tmp_793;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_795 <= _tmp_794;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_796 <= _tmp_795;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_797 <= _tmp_796;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_798 <= _mul_12_sink_busy;
      end 
      if(!_mul_12_sink_busy && _tmp_798) begin
        _mul_12_busy_reg <= 0;
      end 
      if(_mul_12_source_busy) begin
        _mul_12_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_12_fsm_1 = 1;
  localparam _mul_12_fsm_2 = 2;
  localparam _mul_12_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_12_fsm <= _mul_12_fsm_init;
      _mul_12_source_start <= 0;
      _mul_12_source_busy <= 0;
      _mul_12_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_12_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_12_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_12_stream_oready && _tmp_767) begin
        _mul_12_stream_ivalid <= 1;
      end 
      if(_mul_12_stream_oready && 1'd0) begin
        _mul_12_stream_ivalid <= 0;
      end 
      case(_mul_12_fsm)
        _mul_12_fsm_init: begin
          if(_mul_12_run_flag) begin
            _mul_12_source_start <= 1;
          end 
          if(_mul_12_run_flag) begin
            _mul_12_fsm <= _mul_12_fsm_1;
          end 
        end
        _mul_12_fsm_1: begin
          if(_mul_12_source_start && _mul_12_stream_oready) begin
            _mul_12_source_start <= 0;
            _mul_12_source_busy <= 1;
          end 
          if(_mul_12_source_start && _mul_12_stream_oready) begin
            _mul_12_fsm <= _mul_12_fsm_2;
          end 
        end
        _mul_12_fsm_2: begin
          if(_mul_12_stream_oready) begin
            _mul_12_fsm <= _mul_12_fsm_3;
          end 
        end
        _mul_12_fsm_3: begin
          if(_mul_12_stream_oready && 1'd0) begin
            _mul_12_source_busy <= 0;
          end 
          if(_mul_12_stream_oready && 1'd0 && _mul_12_run_flag) begin
            _mul_12_source_start <= 1;
          end 
          if(_mul_12_stream_oready && 1'd0) begin
            _mul_12_fsm <= _mul_12_fsm_init;
          end 
          if(_mul_12_stream_oready && 1'd0 && _mul_12_run_flag) begin
            _mul_12_fsm <= _mul_12_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_13_x_source_ram_renable <= 0;
      _mul_13_x_source_fifo_deq <= 0;
      _mul_13_x_idle <= 1;
      _mul_13_y_source_ram_renable <= 0;
      _mul_13_y_source_fifo_deq <= 0;
      _mul_13_y_idle <= 1;
      _mul_13_rshift_source_ram_renable <= 0;
      _mul_13_rshift_source_fifo_deq <= 0;
      _mul_13_rshift_idle <= 1;
      _mul_13_z_sink_wenable <= 0;
      _mul_13_z_sink_fifo_enq <= 0;
      __mul_13_stream_ivalid_1 <= 0;
      __mul_13_stream_ivalid_2 <= 0;
      __mul_13_stream_ivalid_3 <= 0;
      __mul_13_stream_ivalid_4 <= 0;
      __mul_13_stream_ivalid_5 <= 0;
      __mul_13_stream_ivalid_6 <= 0;
      __mul_13_stream_ivalid_7 <= 0;
      __mul_13_stream_ivalid_8 <= 0;
      _greaterthan_data_244 <= 0;
      _minus_data_246 <= 0;
      _greatereq_data_257 <= 0;
      __delay_data_816__variable_241 <= 0;
      __delay_data_819__variable_242 <= 0;
      __delay_data_822__variable_243 <= 0;
      _sll_data_248 <= 0;
      __delay_data_813_greaterthan_244 <= 0;
      __delay_data_814_greatereq_257 <= 0;
      __delay_data_817__delay_816__variable_241 <= 0;
      __delay_data_820__delay_819__variable_242 <= 0;
      __delay_data_823__delay_822__variable_243 <= 0;
      _cond_data_254 <= 0;
      __delay_data_815__delay_814_greatereq_257 <= 0;
      __delay_data_818__delay_817__delay_816__variable_241 <= 0;
      __delay_data_821__delay_820__delay_819__variable_242 <= 0;
      __delay_data_824__delay_823__delay_822__variable_243 <= 0;
      __muladd_madd_odata_reg_260 <= 0;
      __delay_data_825__delay_824__delay_823____variable_243 <= 0;
      __delay_data_826__delay_825__delay_824____variable_243 <= 0;
      __delay_data_827__delay_826__delay_825____variable_243 <= 0;
      __delay_data_828__delay_827__delay_826____variable_243 <= 0;
      _sra_data_261 <= 0;
      __variable_wdata_241 <= 0;
      __variable_wdata_242 <= 0;
      __variable_wdata_243 <= 0;
      _tmp_799 <= 0;
      _tmp_800 <= 0;
      _tmp_801 <= 0;
      _tmp_802 <= 0;
      _tmp_803 <= 0;
      _tmp_804 <= 0;
      _tmp_805 <= 0;
      _tmp_806 <= 0;
      _tmp_807 <= 0;
      _tmp_808 <= 0;
      _tmp_809 <= 0;
      _tmp_810 <= 0;
      _tmp_811 <= 0;
      _tmp_812 <= 0;
      _tmp_813 <= 0;
      _tmp_814 <= 0;
      _tmp_815 <= 0;
      _tmp_816 <= 0;
      _tmp_817 <= 0;
      _tmp_818 <= 0;
      _tmp_819 <= 0;
      _tmp_820 <= 0;
      _tmp_821 <= 0;
      _tmp_822 <= 0;
      _tmp_823 <= 0;
      _tmp_824 <= 0;
      _tmp_825 <= 0;
      _tmp_826 <= 0;
      _tmp_827 <= 0;
      _tmp_828 <= 0;
      _tmp_829 <= 0;
      _tmp_830 <= 0;
      _tmp_831 <= 0;
      _tmp_832 <= 0;
      _mul_13_busy_reg <= 0;
    end else begin
      if(_mul_13_stream_oready) begin
        _mul_13_x_source_ram_renable <= 0;
        _mul_13_x_source_fifo_deq <= 0;
      end 
      _mul_13_x_idle <= _mul_13_x_idle;
      if(_mul_13_stream_oready) begin
        _mul_13_y_source_ram_renable <= 0;
        _mul_13_y_source_fifo_deq <= 0;
      end 
      _mul_13_y_idle <= _mul_13_y_idle;
      if(_mul_13_stream_oready) begin
        _mul_13_rshift_source_ram_renable <= 0;
        _mul_13_rshift_source_fifo_deq <= 0;
      end 
      _mul_13_rshift_idle <= _mul_13_rshift_idle;
      if(_mul_13_stream_oready) begin
        _mul_13_z_sink_wenable <= 0;
        _mul_13_z_sink_fifo_enq <= 0;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_1 <= _mul_13_stream_ivalid;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_2 <= __mul_13_stream_ivalid_1;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_3 <= __mul_13_stream_ivalid_2;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_4 <= __mul_13_stream_ivalid_3;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_5 <= __mul_13_stream_ivalid_4;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_6 <= __mul_13_stream_ivalid_5;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_7 <= __mul_13_stream_ivalid_6;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_8 <= __mul_13_stream_ivalid_7;
      end 
      if(_mul_13_stream_oready) begin
        _greaterthan_data_244 <= mul_13_rshift_data > 1'sd0;
      end 
      if(_mul_13_stream_oready) begin
        _minus_data_246 <= mul_13_rshift_data - 2'sd1;
      end 
      if(_mul_13_stream_oready) begin
        _greatereq_data_257 <= mul_13_x_data >= 1'sd0;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_816__variable_241 <= mul_13_x_data;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_819__variable_242 <= mul_13_y_data;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_822__variable_243 <= mul_13_rshift_data;
      end 
      if(_mul_13_stream_oready) begin
        _sll_data_248 <= 2'sd1 << _minus_data_246;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_813_greaterthan_244 <= _greaterthan_data_244;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_814_greatereq_257 <= _greatereq_data_257;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_817__delay_816__variable_241 <= __delay_data_816__variable_241;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_820__delay_819__variable_242 <= __delay_data_819__variable_242;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_823__delay_822__variable_243 <= __delay_data_822__variable_243;
      end 
      if(_mul_13_stream_oready) begin
        _cond_data_254 <= (__delay_data_813_greaterthan_244)? _sll_data_248 : 1'sd0;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_815__delay_814_greatereq_257 <= __delay_data_814_greatereq_257;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_818__delay_817__delay_816__variable_241 <= __delay_data_817__delay_816__variable_241;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_821__delay_820__delay_819__variable_242 <= __delay_data_820__delay_819__variable_242;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_824__delay_823__delay_822__variable_243 <= __delay_data_823__delay_822__variable_243;
      end 
      if(_mul_13_stream_oready) begin
        __muladd_madd_odata_reg_260 <= __muladd_madd_odata_260;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_825__delay_824__delay_823____variable_243 <= __delay_data_824__delay_823__delay_822__variable_243;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_826__delay_825__delay_824____variable_243 <= __delay_data_825__delay_824__delay_823____variable_243;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_827__delay_826__delay_825____variable_243 <= __delay_data_826__delay_825__delay_824____variable_243;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_828__delay_827__delay_826____variable_243 <= __delay_data_827__delay_826__delay_825____variable_243;
      end 
      if(_mul_13_stream_oready) begin
        _sra_data_261 <= __muladd_data_260 >>> __delay_data_828__delay_827__delay_826____variable_243;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_241 <= _cond_data_710;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_242 <= __delay_data_1274_reinterpretcast_677;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_243 <= _plus_data_829;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_799 <= _mul_13_source_start;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_800 <= _tmp_799;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_801 <= _tmp_800;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_802 <= _mul_13_source_start;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_803 <= _tmp_802;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_804 <= _tmp_803;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_805 <= _tmp_804;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_806 <= _tmp_805;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_807 <= _tmp_806;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_808 <= _tmp_807;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_809 <= _tmp_808;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_810 <= _tmp_809;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_811 <= _tmp_810;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_812 <= _mul_13_source_stop;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_813 <= _tmp_812;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_814 <= _tmp_813;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_815 <= _tmp_814;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_816 <= _tmp_815;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_817 <= _tmp_816;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_818 <= _tmp_817;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_819 <= _tmp_818;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_820 <= _tmp_819;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_821 <= _tmp_820;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_822 <= _mul_13_source_busy;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_823 <= _tmp_822;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_824 <= _tmp_823;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_825 <= _tmp_824;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_826 <= _tmp_825;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_827 <= _tmp_826;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_828 <= _tmp_827;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_829 <= _tmp_828;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_830 <= _tmp_829;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_831 <= _tmp_830;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_832 <= _mul_13_sink_busy;
      end 
      if(!_mul_13_sink_busy && _tmp_832) begin
        _mul_13_busy_reg <= 0;
      end 
      if(_mul_13_source_busy) begin
        _mul_13_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_13_fsm_1 = 1;
  localparam _mul_13_fsm_2 = 2;
  localparam _mul_13_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_13_fsm <= _mul_13_fsm_init;
      _mul_13_source_start <= 0;
      _mul_13_source_busy <= 0;
      _mul_13_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_13_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_13_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_13_stream_oready && _tmp_801) begin
        _mul_13_stream_ivalid <= 1;
      end 
      if(_mul_13_stream_oready && 1'd0) begin
        _mul_13_stream_ivalid <= 0;
      end 
      case(_mul_13_fsm)
        _mul_13_fsm_init: begin
          if(_mul_13_run_flag) begin
            _mul_13_source_start <= 1;
          end 
          if(_mul_13_run_flag) begin
            _mul_13_fsm <= _mul_13_fsm_1;
          end 
        end
        _mul_13_fsm_1: begin
          if(_mul_13_source_start && _mul_13_stream_oready) begin
            _mul_13_source_start <= 0;
            _mul_13_source_busy <= 1;
          end 
          if(_mul_13_source_start && _mul_13_stream_oready) begin
            _mul_13_fsm <= _mul_13_fsm_2;
          end 
        end
        _mul_13_fsm_2: begin
          if(_mul_13_stream_oready) begin
            _mul_13_fsm <= _mul_13_fsm_3;
          end 
        end
        _mul_13_fsm_3: begin
          if(_mul_13_stream_oready && 1'd0) begin
            _mul_13_source_busy <= 0;
          end 
          if(_mul_13_stream_oready && 1'd0 && _mul_13_run_flag) begin
            _mul_13_source_start <= 1;
          end 
          if(_mul_13_stream_oready && 1'd0) begin
            _mul_13_fsm <= _mul_13_fsm_init;
          end 
          if(_mul_13_stream_oready && 1'd0 && _mul_13_run_flag) begin
            _mul_13_fsm <= _mul_13_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_14_x_source_ram_renable <= 0;
      _mul_14_x_source_fifo_deq <= 0;
      _mul_14_x_idle <= 1;
      _mul_14_y_source_ram_renable <= 0;
      _mul_14_y_source_fifo_deq <= 0;
      _mul_14_y_idle <= 1;
      _mul_14_rshift_source_ram_renable <= 0;
      _mul_14_rshift_source_fifo_deq <= 0;
      _mul_14_rshift_idle <= 1;
      _mul_14_z_sink_wenable <= 0;
      _mul_14_z_sink_fifo_enq <= 0;
      __mul_14_stream_ivalid_1 <= 0;
      __mul_14_stream_ivalid_2 <= 0;
      __mul_14_stream_ivalid_3 <= 0;
      __mul_14_stream_ivalid_4 <= 0;
      __mul_14_stream_ivalid_5 <= 0;
      __mul_14_stream_ivalid_6 <= 0;
      __mul_14_stream_ivalid_7 <= 0;
      __mul_14_stream_ivalid_8 <= 0;
      _greaterthan_data_265 <= 0;
      _minus_data_267 <= 0;
      _greatereq_data_278 <= 0;
      __delay_data_835__variable_262 <= 0;
      __delay_data_838__variable_263 <= 0;
      __delay_data_841__variable_264 <= 0;
      _sll_data_269 <= 0;
      __delay_data_832_greaterthan_265 <= 0;
      __delay_data_833_greatereq_278 <= 0;
      __delay_data_836__delay_835__variable_262 <= 0;
      __delay_data_839__delay_838__variable_263 <= 0;
      __delay_data_842__delay_841__variable_264 <= 0;
      _cond_data_275 <= 0;
      __delay_data_834__delay_833_greatereq_278 <= 0;
      __delay_data_837__delay_836__delay_835__variable_262 <= 0;
      __delay_data_840__delay_839__delay_838__variable_263 <= 0;
      __delay_data_843__delay_842__delay_841__variable_264 <= 0;
      __muladd_madd_odata_reg_281 <= 0;
      __delay_data_844__delay_843__delay_842____variable_264 <= 0;
      __delay_data_845__delay_844__delay_843____variable_264 <= 0;
      __delay_data_846__delay_845__delay_844____variable_264 <= 0;
      __delay_data_847__delay_846__delay_845____variable_264 <= 0;
      _sra_data_282 <= 0;
      __variable_wdata_262 <= 0;
      __variable_wdata_263 <= 0;
      __variable_wdata_264 <= 0;
      _tmp_833 <= 0;
      _tmp_834 <= 0;
      _tmp_835 <= 0;
      _tmp_836 <= 0;
      _tmp_837 <= 0;
      _tmp_838 <= 0;
      _tmp_839 <= 0;
      _tmp_840 <= 0;
      _tmp_841 <= 0;
      _tmp_842 <= 0;
      _tmp_843 <= 0;
      _tmp_844 <= 0;
      _tmp_845 <= 0;
      _tmp_846 <= 0;
      _tmp_847 <= 0;
      _tmp_848 <= 0;
      _tmp_849 <= 0;
      _tmp_850 <= 0;
      _tmp_851 <= 0;
      _tmp_852 <= 0;
      _tmp_853 <= 0;
      _tmp_854 <= 0;
      _tmp_855 <= 0;
      _tmp_856 <= 0;
      _tmp_857 <= 0;
      _tmp_858 <= 0;
      _tmp_859 <= 0;
      _tmp_860 <= 0;
      _tmp_861 <= 0;
      _tmp_862 <= 0;
      _tmp_863 <= 0;
      _tmp_864 <= 0;
      _tmp_865 <= 0;
      _tmp_866 <= 0;
      _mul_14_busy_reg <= 0;
    end else begin
      if(_mul_14_stream_oready) begin
        _mul_14_x_source_ram_renable <= 0;
        _mul_14_x_source_fifo_deq <= 0;
      end 
      _mul_14_x_idle <= _mul_14_x_idle;
      if(_mul_14_stream_oready) begin
        _mul_14_y_source_ram_renable <= 0;
        _mul_14_y_source_fifo_deq <= 0;
      end 
      _mul_14_y_idle <= _mul_14_y_idle;
      if(_mul_14_stream_oready) begin
        _mul_14_rshift_source_ram_renable <= 0;
        _mul_14_rshift_source_fifo_deq <= 0;
      end 
      _mul_14_rshift_idle <= _mul_14_rshift_idle;
      if(_mul_14_stream_oready) begin
        _mul_14_z_sink_wenable <= 0;
        _mul_14_z_sink_fifo_enq <= 0;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_1 <= _mul_14_stream_ivalid;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_2 <= __mul_14_stream_ivalid_1;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_3 <= __mul_14_stream_ivalid_2;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_4 <= __mul_14_stream_ivalid_3;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_5 <= __mul_14_stream_ivalid_4;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_6 <= __mul_14_stream_ivalid_5;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_7 <= __mul_14_stream_ivalid_6;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_8 <= __mul_14_stream_ivalid_7;
      end 
      if(_mul_14_stream_oready) begin
        _greaterthan_data_265 <= mul_14_rshift_data > 1'sd0;
      end 
      if(_mul_14_stream_oready) begin
        _minus_data_267 <= mul_14_rshift_data - 2'sd1;
      end 
      if(_mul_14_stream_oready) begin
        _greatereq_data_278 <= mul_14_x_data >= 1'sd0;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_835__variable_262 <= mul_14_x_data;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_838__variable_263 <= mul_14_y_data;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_841__variable_264 <= mul_14_rshift_data;
      end 
      if(_mul_14_stream_oready) begin
        _sll_data_269 <= 2'sd1 << _minus_data_267;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_832_greaterthan_265 <= _greaterthan_data_265;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_833_greatereq_278 <= _greatereq_data_278;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_836__delay_835__variable_262 <= __delay_data_835__variable_262;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_839__delay_838__variable_263 <= __delay_data_838__variable_263;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_842__delay_841__variable_264 <= __delay_data_841__variable_264;
      end 
      if(_mul_14_stream_oready) begin
        _cond_data_275 <= (__delay_data_832_greaterthan_265)? _sll_data_269 : 1'sd0;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_834__delay_833_greatereq_278 <= __delay_data_833_greatereq_278;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_837__delay_836__delay_835__variable_262 <= __delay_data_836__delay_835__variable_262;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_840__delay_839__delay_838__variable_263 <= __delay_data_839__delay_838__variable_263;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_843__delay_842__delay_841__variable_264 <= __delay_data_842__delay_841__variable_264;
      end 
      if(_mul_14_stream_oready) begin
        __muladd_madd_odata_reg_281 <= __muladd_madd_odata_281;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_844__delay_843__delay_842____variable_264 <= __delay_data_843__delay_842__delay_841__variable_264;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_845__delay_844__delay_843____variable_264 <= __delay_data_844__delay_843__delay_842____variable_264;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_846__delay_845__delay_844____variable_264 <= __delay_data_845__delay_844__delay_843____variable_264;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_847__delay_846__delay_845____variable_264 <= __delay_data_846__delay_845__delay_844____variable_264;
      end 
      if(_mul_14_stream_oready) begin
        _sra_data_282 <= __muladd_data_281 >>> __delay_data_847__delay_846__delay_845____variable_264;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_262 <= _cond_data_712;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_263 <= __delay_data_1276_reinterpretcast_678;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_264 <= _plus_data_848;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_833 <= _mul_14_source_start;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_834 <= _tmp_833;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_835 <= _tmp_834;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_836 <= _mul_14_source_start;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_837 <= _tmp_836;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_838 <= _tmp_837;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_839 <= _tmp_838;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_840 <= _tmp_839;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_841 <= _tmp_840;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_842 <= _tmp_841;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_843 <= _tmp_842;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_844 <= _tmp_843;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_845 <= _tmp_844;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_846 <= _mul_14_source_stop;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_847 <= _tmp_846;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_848 <= _tmp_847;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_849 <= _tmp_848;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_850 <= _tmp_849;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_851 <= _tmp_850;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_852 <= _tmp_851;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_853 <= _tmp_852;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_854 <= _tmp_853;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_855 <= _tmp_854;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_856 <= _mul_14_source_busy;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_857 <= _tmp_856;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_858 <= _tmp_857;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_859 <= _tmp_858;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_860 <= _tmp_859;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_861 <= _tmp_860;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_862 <= _tmp_861;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_863 <= _tmp_862;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_864 <= _tmp_863;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_865 <= _tmp_864;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_866 <= _mul_14_sink_busy;
      end 
      if(!_mul_14_sink_busy && _tmp_866) begin
        _mul_14_busy_reg <= 0;
      end 
      if(_mul_14_source_busy) begin
        _mul_14_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_14_fsm_1 = 1;
  localparam _mul_14_fsm_2 = 2;
  localparam _mul_14_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_14_fsm <= _mul_14_fsm_init;
      _mul_14_source_start <= 0;
      _mul_14_source_busy <= 0;
      _mul_14_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_14_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_14_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_14_stream_oready && _tmp_835) begin
        _mul_14_stream_ivalid <= 1;
      end 
      if(_mul_14_stream_oready && 1'd0) begin
        _mul_14_stream_ivalid <= 0;
      end 
      case(_mul_14_fsm)
        _mul_14_fsm_init: begin
          if(_mul_14_run_flag) begin
            _mul_14_source_start <= 1;
          end 
          if(_mul_14_run_flag) begin
            _mul_14_fsm <= _mul_14_fsm_1;
          end 
        end
        _mul_14_fsm_1: begin
          if(_mul_14_source_start && _mul_14_stream_oready) begin
            _mul_14_source_start <= 0;
            _mul_14_source_busy <= 1;
          end 
          if(_mul_14_source_start && _mul_14_stream_oready) begin
            _mul_14_fsm <= _mul_14_fsm_2;
          end 
        end
        _mul_14_fsm_2: begin
          if(_mul_14_stream_oready) begin
            _mul_14_fsm <= _mul_14_fsm_3;
          end 
        end
        _mul_14_fsm_3: begin
          if(_mul_14_stream_oready && 1'd0) begin
            _mul_14_source_busy <= 0;
          end 
          if(_mul_14_stream_oready && 1'd0 && _mul_14_run_flag) begin
            _mul_14_source_start <= 1;
          end 
          if(_mul_14_stream_oready && 1'd0) begin
            _mul_14_fsm <= _mul_14_fsm_init;
          end 
          if(_mul_14_stream_oready && 1'd0 && _mul_14_run_flag) begin
            _mul_14_fsm <= _mul_14_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_15_x_source_ram_renable <= 0;
      _mul_15_x_source_fifo_deq <= 0;
      _mul_15_x_idle <= 1;
      _mul_15_y_source_ram_renable <= 0;
      _mul_15_y_source_fifo_deq <= 0;
      _mul_15_y_idle <= 1;
      _mul_15_rshift_source_ram_renable <= 0;
      _mul_15_rshift_source_fifo_deq <= 0;
      _mul_15_rshift_idle <= 1;
      _mul_15_z_sink_wenable <= 0;
      _mul_15_z_sink_fifo_enq <= 0;
      __mul_15_stream_ivalid_1 <= 0;
      __mul_15_stream_ivalid_2 <= 0;
      __mul_15_stream_ivalid_3 <= 0;
      __mul_15_stream_ivalid_4 <= 0;
      __mul_15_stream_ivalid_5 <= 0;
      __mul_15_stream_ivalid_6 <= 0;
      __mul_15_stream_ivalid_7 <= 0;
      __mul_15_stream_ivalid_8 <= 0;
      _greaterthan_data_286 <= 0;
      _minus_data_288 <= 0;
      _greatereq_data_299 <= 0;
      __delay_data_854__variable_283 <= 0;
      __delay_data_857__variable_284 <= 0;
      __delay_data_860__variable_285 <= 0;
      _sll_data_290 <= 0;
      __delay_data_851_greaterthan_286 <= 0;
      __delay_data_852_greatereq_299 <= 0;
      __delay_data_855__delay_854__variable_283 <= 0;
      __delay_data_858__delay_857__variable_284 <= 0;
      __delay_data_861__delay_860__variable_285 <= 0;
      _cond_data_296 <= 0;
      __delay_data_853__delay_852_greatereq_299 <= 0;
      __delay_data_856__delay_855__delay_854__variable_283 <= 0;
      __delay_data_859__delay_858__delay_857__variable_284 <= 0;
      __delay_data_862__delay_861__delay_860__variable_285 <= 0;
      __muladd_madd_odata_reg_302 <= 0;
      __delay_data_863__delay_862__delay_861____variable_285 <= 0;
      __delay_data_864__delay_863__delay_862____variable_285 <= 0;
      __delay_data_865__delay_864__delay_863____variable_285 <= 0;
      __delay_data_866__delay_865__delay_864____variable_285 <= 0;
      _sra_data_303 <= 0;
      __variable_wdata_283 <= 0;
      __variable_wdata_284 <= 0;
      __variable_wdata_285 <= 0;
      _tmp_867 <= 0;
      _tmp_868 <= 0;
      _tmp_869 <= 0;
      _tmp_870 <= 0;
      _tmp_871 <= 0;
      _tmp_872 <= 0;
      _tmp_873 <= 0;
      _tmp_874 <= 0;
      _tmp_875 <= 0;
      _tmp_876 <= 0;
      _tmp_877 <= 0;
      _tmp_878 <= 0;
      _tmp_879 <= 0;
      _tmp_880 <= 0;
      _tmp_881 <= 0;
      _tmp_882 <= 0;
      _tmp_883 <= 0;
      _tmp_884 <= 0;
      _tmp_885 <= 0;
      _tmp_886 <= 0;
      _tmp_887 <= 0;
      _tmp_888 <= 0;
      _tmp_889 <= 0;
      _tmp_890 <= 0;
      _tmp_891 <= 0;
      _tmp_892 <= 0;
      _tmp_893 <= 0;
      _tmp_894 <= 0;
      _tmp_895 <= 0;
      _tmp_896 <= 0;
      _tmp_897 <= 0;
      _tmp_898 <= 0;
      _tmp_899 <= 0;
      _tmp_900 <= 0;
      _mul_15_busy_reg <= 0;
    end else begin
      if(_mul_15_stream_oready) begin
        _mul_15_x_source_ram_renable <= 0;
        _mul_15_x_source_fifo_deq <= 0;
      end 
      _mul_15_x_idle <= _mul_15_x_idle;
      if(_mul_15_stream_oready) begin
        _mul_15_y_source_ram_renable <= 0;
        _mul_15_y_source_fifo_deq <= 0;
      end 
      _mul_15_y_idle <= _mul_15_y_idle;
      if(_mul_15_stream_oready) begin
        _mul_15_rshift_source_ram_renable <= 0;
        _mul_15_rshift_source_fifo_deq <= 0;
      end 
      _mul_15_rshift_idle <= _mul_15_rshift_idle;
      if(_mul_15_stream_oready) begin
        _mul_15_z_sink_wenable <= 0;
        _mul_15_z_sink_fifo_enq <= 0;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_1 <= _mul_15_stream_ivalid;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_2 <= __mul_15_stream_ivalid_1;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_3 <= __mul_15_stream_ivalid_2;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_4 <= __mul_15_stream_ivalid_3;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_5 <= __mul_15_stream_ivalid_4;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_6 <= __mul_15_stream_ivalid_5;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_7 <= __mul_15_stream_ivalid_6;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_8 <= __mul_15_stream_ivalid_7;
      end 
      if(_mul_15_stream_oready) begin
        _greaterthan_data_286 <= mul_15_rshift_data > 1'sd0;
      end 
      if(_mul_15_stream_oready) begin
        _minus_data_288 <= mul_15_rshift_data - 2'sd1;
      end 
      if(_mul_15_stream_oready) begin
        _greatereq_data_299 <= mul_15_x_data >= 1'sd0;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_854__variable_283 <= mul_15_x_data;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_857__variable_284 <= mul_15_y_data;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_860__variable_285 <= mul_15_rshift_data;
      end 
      if(_mul_15_stream_oready) begin
        _sll_data_290 <= 2'sd1 << _minus_data_288;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_851_greaterthan_286 <= _greaterthan_data_286;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_852_greatereq_299 <= _greatereq_data_299;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_855__delay_854__variable_283 <= __delay_data_854__variable_283;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_858__delay_857__variable_284 <= __delay_data_857__variable_284;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_861__delay_860__variable_285 <= __delay_data_860__variable_285;
      end 
      if(_mul_15_stream_oready) begin
        _cond_data_296 <= (__delay_data_851_greaterthan_286)? _sll_data_290 : 1'sd0;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_853__delay_852_greatereq_299 <= __delay_data_852_greatereq_299;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_856__delay_855__delay_854__variable_283 <= __delay_data_855__delay_854__variable_283;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_859__delay_858__delay_857__variable_284 <= __delay_data_858__delay_857__variable_284;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_862__delay_861__delay_860__variable_285 <= __delay_data_861__delay_860__variable_285;
      end 
      if(_mul_15_stream_oready) begin
        __muladd_madd_odata_reg_302 <= __muladd_madd_odata_302;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_863__delay_862__delay_861____variable_285 <= __delay_data_862__delay_861__delay_860__variable_285;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_864__delay_863__delay_862____variable_285 <= __delay_data_863__delay_862__delay_861____variable_285;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_865__delay_864__delay_863____variable_285 <= __delay_data_864__delay_863__delay_862____variable_285;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_866__delay_865__delay_864____variable_285 <= __delay_data_865__delay_864__delay_863____variable_285;
      end 
      if(_mul_15_stream_oready) begin
        _sra_data_303 <= __muladd_data_302 >>> __delay_data_866__delay_865__delay_864____variable_285;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_283 <= _cond_data_714;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_284 <= __delay_data_1278_reinterpretcast_679;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_285 <= _plus_data_867;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_867 <= _mul_15_source_start;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_868 <= _tmp_867;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_869 <= _tmp_868;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_870 <= _mul_15_source_start;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_871 <= _tmp_870;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_872 <= _tmp_871;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_873 <= _tmp_872;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_874 <= _tmp_873;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_875 <= _tmp_874;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_876 <= _tmp_875;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_877 <= _tmp_876;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_878 <= _tmp_877;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_879 <= _tmp_878;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_880 <= _mul_15_source_stop;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_881 <= _tmp_880;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_882 <= _tmp_881;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_883 <= _tmp_882;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_884 <= _tmp_883;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_885 <= _tmp_884;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_886 <= _tmp_885;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_887 <= _tmp_886;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_888 <= _tmp_887;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_889 <= _tmp_888;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_890 <= _mul_15_source_busy;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_891 <= _tmp_890;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_892 <= _tmp_891;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_893 <= _tmp_892;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_894 <= _tmp_893;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_895 <= _tmp_894;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_896 <= _tmp_895;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_897 <= _tmp_896;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_898 <= _tmp_897;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_899 <= _tmp_898;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_900 <= _mul_15_sink_busy;
      end 
      if(!_mul_15_sink_busy && _tmp_900) begin
        _mul_15_busy_reg <= 0;
      end 
      if(_mul_15_source_busy) begin
        _mul_15_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_15_fsm_1 = 1;
  localparam _mul_15_fsm_2 = 2;
  localparam _mul_15_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_15_fsm <= _mul_15_fsm_init;
      _mul_15_source_start <= 0;
      _mul_15_source_busy <= 0;
      _mul_15_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_15_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_15_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_15_stream_oready && _tmp_869) begin
        _mul_15_stream_ivalid <= 1;
      end 
      if(_mul_15_stream_oready && 1'd0) begin
        _mul_15_stream_ivalid <= 0;
      end 
      case(_mul_15_fsm)
        _mul_15_fsm_init: begin
          if(_mul_15_run_flag) begin
            _mul_15_source_start <= 1;
          end 
          if(_mul_15_run_flag) begin
            _mul_15_fsm <= _mul_15_fsm_1;
          end 
        end
        _mul_15_fsm_1: begin
          if(_mul_15_source_start && _mul_15_stream_oready) begin
            _mul_15_source_start <= 0;
            _mul_15_source_busy <= 1;
          end 
          if(_mul_15_source_start && _mul_15_stream_oready) begin
            _mul_15_fsm <= _mul_15_fsm_2;
          end 
        end
        _mul_15_fsm_2: begin
          if(_mul_15_stream_oready) begin
            _mul_15_fsm <= _mul_15_fsm_3;
          end 
        end
        _mul_15_fsm_3: begin
          if(_mul_15_stream_oready && 1'd0) begin
            _mul_15_source_busy <= 0;
          end 
          if(_mul_15_stream_oready && 1'd0 && _mul_15_run_flag) begin
            _mul_15_source_start <= 1;
          end 
          if(_mul_15_stream_oready && 1'd0) begin
            _mul_15_fsm <= _mul_15_fsm_init;
          end 
          if(_mul_15_stream_oready && 1'd0 && _mul_15_run_flag) begin
            _mul_15_fsm <= _mul_15_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_16_x_source_ram_renable <= 0;
      _mul_16_x_source_fifo_deq <= 0;
      _mul_16_x_idle <= 1;
      _mul_16_y_source_ram_renable <= 0;
      _mul_16_y_source_fifo_deq <= 0;
      _mul_16_y_idle <= 1;
      _mul_16_rshift_source_ram_renable <= 0;
      _mul_16_rshift_source_fifo_deq <= 0;
      _mul_16_rshift_idle <= 1;
      _mul_16_z_sink_wenable <= 0;
      _mul_16_z_sink_fifo_enq <= 0;
      __mul_16_stream_ivalid_1 <= 0;
      __mul_16_stream_ivalid_2 <= 0;
      __mul_16_stream_ivalid_3 <= 0;
      __mul_16_stream_ivalid_4 <= 0;
      __mul_16_stream_ivalid_5 <= 0;
      __mul_16_stream_ivalid_6 <= 0;
      __mul_16_stream_ivalid_7 <= 0;
      __mul_16_stream_ivalid_8 <= 0;
      _greaterthan_data_307 <= 0;
      _minus_data_309 <= 0;
      _greatereq_data_320 <= 0;
      __delay_data_873__variable_304 <= 0;
      __delay_data_876__variable_305 <= 0;
      __delay_data_879__variable_306 <= 0;
      _sll_data_311 <= 0;
      __delay_data_870_greaterthan_307 <= 0;
      __delay_data_871_greatereq_320 <= 0;
      __delay_data_874__delay_873__variable_304 <= 0;
      __delay_data_877__delay_876__variable_305 <= 0;
      __delay_data_880__delay_879__variable_306 <= 0;
      _cond_data_317 <= 0;
      __delay_data_872__delay_871_greatereq_320 <= 0;
      __delay_data_875__delay_874__delay_873__variable_304 <= 0;
      __delay_data_878__delay_877__delay_876__variable_305 <= 0;
      __delay_data_881__delay_880__delay_879__variable_306 <= 0;
      __muladd_madd_odata_reg_323 <= 0;
      __delay_data_882__delay_881__delay_880____variable_306 <= 0;
      __delay_data_883__delay_882__delay_881____variable_306 <= 0;
      __delay_data_884__delay_883__delay_882____variable_306 <= 0;
      __delay_data_885__delay_884__delay_883____variable_306 <= 0;
      _sra_data_324 <= 0;
      __variable_wdata_304 <= 0;
      __variable_wdata_305 <= 0;
      __variable_wdata_306 <= 0;
      _tmp_901 <= 0;
      _tmp_902 <= 0;
      _tmp_903 <= 0;
      _tmp_904 <= 0;
      _tmp_905 <= 0;
      _tmp_906 <= 0;
      _tmp_907 <= 0;
      _tmp_908 <= 0;
      _tmp_909 <= 0;
      _tmp_910 <= 0;
      _tmp_911 <= 0;
      _tmp_912 <= 0;
      _tmp_913 <= 0;
      _tmp_914 <= 0;
      _tmp_915 <= 0;
      _tmp_916 <= 0;
      _tmp_917 <= 0;
      _tmp_918 <= 0;
      _tmp_919 <= 0;
      _tmp_920 <= 0;
      _tmp_921 <= 0;
      _tmp_922 <= 0;
      _tmp_923 <= 0;
      _tmp_924 <= 0;
      _tmp_925 <= 0;
      _tmp_926 <= 0;
      _tmp_927 <= 0;
      _tmp_928 <= 0;
      _tmp_929 <= 0;
      _tmp_930 <= 0;
      _tmp_931 <= 0;
      _tmp_932 <= 0;
      _tmp_933 <= 0;
      _tmp_934 <= 0;
      _mul_16_busy_reg <= 0;
    end else begin
      if(_mul_16_stream_oready) begin
        _mul_16_x_source_ram_renable <= 0;
        _mul_16_x_source_fifo_deq <= 0;
      end 
      _mul_16_x_idle <= _mul_16_x_idle;
      if(_mul_16_stream_oready) begin
        _mul_16_y_source_ram_renable <= 0;
        _mul_16_y_source_fifo_deq <= 0;
      end 
      _mul_16_y_idle <= _mul_16_y_idle;
      if(_mul_16_stream_oready) begin
        _mul_16_rshift_source_ram_renable <= 0;
        _mul_16_rshift_source_fifo_deq <= 0;
      end 
      _mul_16_rshift_idle <= _mul_16_rshift_idle;
      if(_mul_16_stream_oready) begin
        _mul_16_z_sink_wenable <= 0;
        _mul_16_z_sink_fifo_enq <= 0;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_1 <= _mul_16_stream_ivalid;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_2 <= __mul_16_stream_ivalid_1;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_3 <= __mul_16_stream_ivalid_2;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_4 <= __mul_16_stream_ivalid_3;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_5 <= __mul_16_stream_ivalid_4;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_6 <= __mul_16_stream_ivalid_5;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_7 <= __mul_16_stream_ivalid_6;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_8 <= __mul_16_stream_ivalid_7;
      end 
      if(_mul_16_stream_oready) begin
        _greaterthan_data_307 <= mul_16_rshift_data > 1'sd0;
      end 
      if(_mul_16_stream_oready) begin
        _minus_data_309 <= mul_16_rshift_data - 2'sd1;
      end 
      if(_mul_16_stream_oready) begin
        _greatereq_data_320 <= mul_16_x_data >= 1'sd0;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_873__variable_304 <= mul_16_x_data;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_876__variable_305 <= mul_16_y_data;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_879__variable_306 <= mul_16_rshift_data;
      end 
      if(_mul_16_stream_oready) begin
        _sll_data_311 <= 2'sd1 << _minus_data_309;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_870_greaterthan_307 <= _greaterthan_data_307;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_871_greatereq_320 <= _greatereq_data_320;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_874__delay_873__variable_304 <= __delay_data_873__variable_304;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_877__delay_876__variable_305 <= __delay_data_876__variable_305;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_880__delay_879__variable_306 <= __delay_data_879__variable_306;
      end 
      if(_mul_16_stream_oready) begin
        _cond_data_317 <= (__delay_data_870_greaterthan_307)? _sll_data_311 : 1'sd0;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_872__delay_871_greatereq_320 <= __delay_data_871_greatereq_320;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_875__delay_874__delay_873__variable_304 <= __delay_data_874__delay_873__variable_304;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_878__delay_877__delay_876__variable_305 <= __delay_data_877__delay_876__variable_305;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_881__delay_880__delay_879__variable_306 <= __delay_data_880__delay_879__variable_306;
      end 
      if(_mul_16_stream_oready) begin
        __muladd_madd_odata_reg_323 <= __muladd_madd_odata_323;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_882__delay_881__delay_880____variable_306 <= __delay_data_881__delay_880__delay_879__variable_306;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_883__delay_882__delay_881____variable_306 <= __delay_data_882__delay_881__delay_880____variable_306;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_884__delay_883__delay_882____variable_306 <= __delay_data_883__delay_882__delay_881____variable_306;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_885__delay_884__delay_883____variable_306 <= __delay_data_884__delay_883__delay_882____variable_306;
      end 
      if(_mul_16_stream_oready) begin
        _sra_data_324 <= __muladd_data_323 >>> __delay_data_885__delay_884__delay_883____variable_306;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_304 <= _cond_data_716;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_305 <= __delay_data_1280_reinterpretcast_680;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_306 <= _plus_data_886;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_901 <= _mul_16_source_start;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_902 <= _tmp_901;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_903 <= _tmp_902;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_904 <= _mul_16_source_start;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_905 <= _tmp_904;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_906 <= _tmp_905;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_907 <= _tmp_906;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_908 <= _tmp_907;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_909 <= _tmp_908;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_910 <= _tmp_909;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_911 <= _tmp_910;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_912 <= _tmp_911;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_913 <= _tmp_912;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_914 <= _mul_16_source_stop;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_915 <= _tmp_914;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_916 <= _tmp_915;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_917 <= _tmp_916;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_918 <= _tmp_917;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_919 <= _tmp_918;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_920 <= _tmp_919;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_921 <= _tmp_920;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_922 <= _tmp_921;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_923 <= _tmp_922;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_924 <= _mul_16_source_busy;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_925 <= _tmp_924;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_926 <= _tmp_925;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_927 <= _tmp_926;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_928 <= _tmp_927;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_929 <= _tmp_928;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_930 <= _tmp_929;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_931 <= _tmp_930;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_932 <= _tmp_931;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_933 <= _tmp_932;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_934 <= _mul_16_sink_busy;
      end 
      if(!_mul_16_sink_busy && _tmp_934) begin
        _mul_16_busy_reg <= 0;
      end 
      if(_mul_16_source_busy) begin
        _mul_16_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_16_fsm_1 = 1;
  localparam _mul_16_fsm_2 = 2;
  localparam _mul_16_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_16_fsm <= _mul_16_fsm_init;
      _mul_16_source_start <= 0;
      _mul_16_source_busy <= 0;
      _mul_16_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_16_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_16_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_16_stream_oready && _tmp_903) begin
        _mul_16_stream_ivalid <= 1;
      end 
      if(_mul_16_stream_oready && 1'd0) begin
        _mul_16_stream_ivalid <= 0;
      end 
      case(_mul_16_fsm)
        _mul_16_fsm_init: begin
          if(_mul_16_run_flag) begin
            _mul_16_source_start <= 1;
          end 
          if(_mul_16_run_flag) begin
            _mul_16_fsm <= _mul_16_fsm_1;
          end 
        end
        _mul_16_fsm_1: begin
          if(_mul_16_source_start && _mul_16_stream_oready) begin
            _mul_16_source_start <= 0;
            _mul_16_source_busy <= 1;
          end 
          if(_mul_16_source_start && _mul_16_stream_oready) begin
            _mul_16_fsm <= _mul_16_fsm_2;
          end 
        end
        _mul_16_fsm_2: begin
          if(_mul_16_stream_oready) begin
            _mul_16_fsm <= _mul_16_fsm_3;
          end 
        end
        _mul_16_fsm_3: begin
          if(_mul_16_stream_oready && 1'd0) begin
            _mul_16_source_busy <= 0;
          end 
          if(_mul_16_stream_oready && 1'd0 && _mul_16_run_flag) begin
            _mul_16_source_start <= 1;
          end 
          if(_mul_16_stream_oready && 1'd0) begin
            _mul_16_fsm <= _mul_16_fsm_init;
          end 
          if(_mul_16_stream_oready && 1'd0 && _mul_16_run_flag) begin
            _mul_16_fsm <= _mul_16_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_17_x_source_ram_renable <= 0;
      __reduce_max_17_x_source_fifo_deq <= 0;
      __reduce_max_17_x_idle <= 1;
      __reduce_max_17_data_sink_wenable <= 0;
      __reduce_max_17_data_sink_fifo_enq <= 0;
      __reduce_max_17_valid_sink_wenable <= 0;
      __reduce_max_17_valid_sink_fifo_enq <= 0;
      ___reduce_max_17_stream_ivalid_1 <= 0;
      _reducemax_data_328 <= -17'sd32768;
      _reducemax_count_328 <= 0;
      _reducemax_prev_count_max_328 <= 0;
      _pulse_data_330 <= 1'sd0;
      _pulse_count_330 <= 0;
      _pulse_prev_count_max_330 <= 0;
      __variable_wdata_327 <= 0;
      __variable_wdata_325 <= 0;
      __variable_wdata_326 <= 0;
      _tmp_1218 <= 0;
      _tmp_1219 <= 0;
      _tmp_1220 <= 0;
      _tmp_1221 <= 0;
      _tmp_1222 <= 0;
      _tmp_1223 <= 0;
      _tmp_1224 <= 0;
      _tmp_1225 <= 0;
      _tmp_1226 <= 0;
      _tmp_1227 <= 0;
      _tmp_1228 <= 0;
      _tmp_1229 <= 0;
      _tmp_1230 <= 0;
      _tmp_1231 <= 0;
      _tmp_1232 <= 0;
      _tmp_1233 <= 0;
      _tmp_1234 <= 0;
      _tmp_1235 <= 0;
      _tmp_1236 <= 0;
      _tmp_1237 <= 0;
      __reduce_max_17_busy_reg <= 0;
    end else begin
      if(__reduce_max_17_stream_oready) begin
        __reduce_max_17_x_source_ram_renable <= 0;
        __reduce_max_17_x_source_fifo_deq <= 0;
      end 
      __reduce_max_17_x_idle <= __reduce_max_17_x_idle;
      if(__reduce_max_17_stream_oready) begin
        __reduce_max_17_data_sink_wenable <= 0;
        __reduce_max_17_data_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_17_stream_oready) begin
        __reduce_max_17_valid_sink_wenable <= 0;
        __reduce_max_17_valid_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_17_stream_oready) begin
        ___reduce_max_17_stream_ivalid_1 <= __reduce_max_17_stream_ivalid;
      end 
      if(__reduce_max_17_stream_ivalid && __reduce_max_17_stream_oready && _reducemax_reset_cond_328) begin
        _reducemax_data_328 <= -17'sd32768;
      end 
      if(__reduce_max_17_stream_ivalid && __reduce_max_17_stream_oready) begin
        _reducemax_count_328 <= (_reducemax_current_count_328 >= _reduce_max_17_size_data - 1)? 0 : _reducemax_current_count_328 + 1;
      end 
      if(__reduce_max_17_stream_ivalid && __reduce_max_17_stream_oready) begin
        _reducemax_prev_count_max_328 <= _reducemax_current_count_328 >= _reduce_max_17_size_data - 1;
      end 
      if(__reduce_max_17_stream_ivalid && __reduce_max_17_stream_oready) begin
        _reducemax_data_328 <= (_reducemax_current_data_328 < _reduce_max_17_x_data)? _reduce_max_17_x_data : _reducemax_current_data_328;
      end 
      if(__reduce_max_17_stream_ivalid && __reduce_max_17_stream_oready && _pulse_reset_cond_330) begin
        _pulse_data_330 <= 1'sd0;
      end 
      if(__reduce_max_17_stream_ivalid && __reduce_max_17_stream_oready) begin
        _pulse_count_330 <= (_pulse_current_count_330 >= _reduce_max_17_size_data - 1)? 0 : _pulse_current_count_330 + 1;
      end 
      if(__reduce_max_17_stream_ivalid && __reduce_max_17_stream_oready) begin
        _pulse_prev_count_max_330 <= _pulse_current_count_330 >= _reduce_max_17_size_data - 1;
      end 
      if(__reduce_max_17_stream_ivalid && __reduce_max_17_stream_oready) begin
        _pulse_data_330 <= _pulse_current_count_330 >= _reduce_max_17_size_data - 1;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_327 <= __delay_data_1395__delay_1394__delay_1393__variable_931;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_325 <= _cond_data_945;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_326 <= __delay_data_1398__delay_1397__delay_1396__variable_928;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1218 <= __reduce_max_17_source_start;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1219 <= _tmp_1218;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1220 <= _tmp_1219;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1221 <= __reduce_max_17_source_start;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1222 <= _tmp_1221;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1223 <= _tmp_1222;
      end 
      if(__reduce_max_17_stream_oready && _tmp_1223) begin
        __variable_wdata_327 <= 1;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1224 <= __reduce_max_17_source_start;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1225 <= _tmp_1224;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1226 <= _tmp_1225;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1227 <= _tmp_1226;
      end 
      if(__reduce_max_17_stream_oready && _tmp_1227) begin
        __variable_wdata_327 <= 0;
      end 
      if(__reduce_max_17_stream_oready && 1'd0) begin
        __variable_wdata_327 <= 1;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1228 <= __reduce_max_17_source_start;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1229 <= _tmp_1228;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1230 <= _tmp_1229;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1231 <= __reduce_max_17_source_stop;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1232 <= _tmp_1231;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1233 <= _tmp_1232;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1234 <= __reduce_max_17_source_busy;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1235 <= _tmp_1234;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1236 <= _tmp_1235;
      end 
      if(__reduce_max_17_stream_oready) begin
        _tmp_1237 <= __reduce_max_17_sink_busy;
      end 
      if(!__reduce_max_17_sink_busy && _tmp_1237) begin
        __reduce_max_17_busy_reg <= 0;
      end 
      if(__reduce_max_17_source_busy) begin
        __reduce_max_17_busy_reg <= 1;
      end 
    end
  end

  localparam __reduce_max_17_fsm_1 = 1;
  localparam __reduce_max_17_fsm_2 = 2;
  localparam __reduce_max_17_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_17_fsm <= __reduce_max_17_fsm_init;
      __reduce_max_17_source_start <= 0;
      __reduce_max_17_source_busy <= 0;
      __reduce_max_17_stream_ivalid <= 0;
    end else begin
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __reduce_max_17_stream_ivalid <= 1'd1;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_busy) begin
        __reduce_max_17_source_busy <= _stream_max_pool_serial_6_source_busy;
      end 
      if(__reduce_max_17_stream_oready && _tmp_1220) begin
        __reduce_max_17_stream_ivalid <= 1;
      end 
      if(__reduce_max_17_stream_oready && 1'd0) begin
        __reduce_max_17_stream_ivalid <= 0;
      end 
      case(__reduce_max_17_fsm)
        __reduce_max_17_fsm_init: begin
          if(__reduce_max_17_run_flag) begin
            __reduce_max_17_source_start <= 1;
          end 
          if(__reduce_max_17_run_flag) begin
            __reduce_max_17_fsm <= __reduce_max_17_fsm_1;
          end 
        end
        __reduce_max_17_fsm_1: begin
          if(__reduce_max_17_source_start && __reduce_max_17_stream_oready) begin
            __reduce_max_17_source_start <= 0;
            __reduce_max_17_source_busy <= 1;
          end 
          if(__reduce_max_17_source_start && __reduce_max_17_stream_oready) begin
            __reduce_max_17_fsm <= __reduce_max_17_fsm_2;
          end 
        end
        __reduce_max_17_fsm_2: begin
          if(__reduce_max_17_stream_oready) begin
            __reduce_max_17_fsm <= __reduce_max_17_fsm_3;
          end 
        end
        __reduce_max_17_fsm_3: begin
          if(__reduce_max_17_stream_oready && 1'd0) begin
            __reduce_max_17_source_busy <= 0;
          end 
          if(__reduce_max_17_stream_oready && 1'd0 && __reduce_max_17_run_flag) begin
            __reduce_max_17_source_start <= 1;
          end 
          if(__reduce_max_17_stream_oready && 1'd0) begin
            __reduce_max_17_fsm <= __reduce_max_17_fsm_init;
          end 
          if(__reduce_max_17_stream_oready && 1'd0 && __reduce_max_17_run_flag) begin
            __reduce_max_17_fsm <= __reduce_max_17_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_18_x_source_ram_renable <= 0;
      __reduce_max_18_x_source_fifo_deq <= 0;
      __reduce_max_18_x_idle <= 1;
      __reduce_max_18_data_sink_wenable <= 0;
      __reduce_max_18_data_sink_fifo_enq <= 0;
      __reduce_max_18_valid_sink_wenable <= 0;
      __reduce_max_18_valid_sink_fifo_enq <= 0;
      ___reduce_max_18_stream_ivalid_1 <= 0;
      _reducemax_data_335 <= -17'sd32768;
      _reducemax_count_335 <= 0;
      _reducemax_prev_count_max_335 <= 0;
      _pulse_data_337 <= 1'sd0;
      _pulse_count_337 <= 0;
      _pulse_prev_count_max_337 <= 0;
      __variable_wdata_334 <= 0;
      __variable_wdata_332 <= 0;
      __variable_wdata_333 <= 0;
      _tmp_1238 <= 0;
      _tmp_1239 <= 0;
      _tmp_1240 <= 0;
      _tmp_1241 <= 0;
      _tmp_1242 <= 0;
      _tmp_1243 <= 0;
      _tmp_1244 <= 0;
      _tmp_1245 <= 0;
      _tmp_1246 <= 0;
      _tmp_1247 <= 0;
      _tmp_1248 <= 0;
      _tmp_1249 <= 0;
      _tmp_1250 <= 0;
      _tmp_1251 <= 0;
      _tmp_1252 <= 0;
      _tmp_1253 <= 0;
      _tmp_1254 <= 0;
      _tmp_1255 <= 0;
      _tmp_1256 <= 0;
      _tmp_1257 <= 0;
      __reduce_max_18_busy_reg <= 0;
    end else begin
      if(__reduce_max_18_stream_oready) begin
        __reduce_max_18_x_source_ram_renable <= 0;
        __reduce_max_18_x_source_fifo_deq <= 0;
      end 
      __reduce_max_18_x_idle <= __reduce_max_18_x_idle;
      if(__reduce_max_18_stream_oready) begin
        __reduce_max_18_data_sink_wenable <= 0;
        __reduce_max_18_data_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_18_stream_oready) begin
        __reduce_max_18_valid_sink_wenable <= 0;
        __reduce_max_18_valid_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_18_stream_oready) begin
        ___reduce_max_18_stream_ivalid_1 <= __reduce_max_18_stream_ivalid;
      end 
      if(__reduce_max_18_stream_ivalid && __reduce_max_18_stream_oready && _reducemax_reset_cond_335) begin
        _reducemax_data_335 <= -17'sd32768;
      end 
      if(__reduce_max_18_stream_ivalid && __reduce_max_18_stream_oready) begin
        _reducemax_count_335 <= (_reducemax_current_count_335 >= _reduce_max_18_size_data - 1)? 0 : _reducemax_current_count_335 + 1;
      end 
      if(__reduce_max_18_stream_ivalid && __reduce_max_18_stream_oready) begin
        _reducemax_prev_count_max_335 <= _reducemax_current_count_335 >= _reduce_max_18_size_data - 1;
      end 
      if(__reduce_max_18_stream_ivalid && __reduce_max_18_stream_oready) begin
        _reducemax_data_335 <= (_reducemax_current_data_335 < _reduce_max_18_x_data)? _reduce_max_18_x_data : _reducemax_current_data_335;
      end 
      if(__reduce_max_18_stream_ivalid && __reduce_max_18_stream_oready && _pulse_reset_cond_337) begin
        _pulse_data_337 <= 1'sd0;
      end 
      if(__reduce_max_18_stream_ivalid && __reduce_max_18_stream_oready) begin
        _pulse_count_337 <= (_pulse_current_count_337 >= _reduce_max_18_size_data - 1)? 0 : _pulse_current_count_337 + 1;
      end 
      if(__reduce_max_18_stream_ivalid && __reduce_max_18_stream_oready) begin
        _pulse_prev_count_max_337 <= _pulse_current_count_337 >= _reduce_max_18_size_data - 1;
      end 
      if(__reduce_max_18_stream_ivalid && __reduce_max_18_stream_oready) begin
        _pulse_data_337 <= _pulse_current_count_337 >= _reduce_max_18_size_data - 1;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_334 <= __delay_data_1395__delay_1394__delay_1393__variable_931;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_332 <= _cond_data_950;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_333 <= __delay_data_1398__delay_1397__delay_1396__variable_928;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1238 <= __reduce_max_18_source_start;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1239 <= _tmp_1238;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1240 <= _tmp_1239;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1241 <= __reduce_max_18_source_start;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1242 <= _tmp_1241;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1243 <= _tmp_1242;
      end 
      if(__reduce_max_18_stream_oready && _tmp_1243) begin
        __variable_wdata_334 <= 1;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1244 <= __reduce_max_18_source_start;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1245 <= _tmp_1244;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1246 <= _tmp_1245;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1247 <= _tmp_1246;
      end 
      if(__reduce_max_18_stream_oready && _tmp_1247) begin
        __variable_wdata_334 <= 0;
      end 
      if(__reduce_max_18_stream_oready && 1'd0) begin
        __variable_wdata_334 <= 1;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1248 <= __reduce_max_18_source_start;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1249 <= _tmp_1248;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1250 <= _tmp_1249;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1251 <= __reduce_max_18_source_stop;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1252 <= _tmp_1251;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1253 <= _tmp_1252;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1254 <= __reduce_max_18_source_busy;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1255 <= _tmp_1254;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1256 <= _tmp_1255;
      end 
      if(__reduce_max_18_stream_oready) begin
        _tmp_1257 <= __reduce_max_18_sink_busy;
      end 
      if(!__reduce_max_18_sink_busy && _tmp_1257) begin
        __reduce_max_18_busy_reg <= 0;
      end 
      if(__reduce_max_18_source_busy) begin
        __reduce_max_18_busy_reg <= 1;
      end 
    end
  end

  localparam __reduce_max_18_fsm_1 = 1;
  localparam __reduce_max_18_fsm_2 = 2;
  localparam __reduce_max_18_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_18_fsm <= __reduce_max_18_fsm_init;
      __reduce_max_18_source_start <= 0;
      __reduce_max_18_source_busy <= 0;
      __reduce_max_18_stream_ivalid <= 0;
    end else begin
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __reduce_max_18_stream_ivalid <= 1'd1;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_busy) begin
        __reduce_max_18_source_busy <= _stream_max_pool_serial_6_source_busy;
      end 
      if(__reduce_max_18_stream_oready && _tmp_1240) begin
        __reduce_max_18_stream_ivalid <= 1;
      end 
      if(__reduce_max_18_stream_oready && 1'd0) begin
        __reduce_max_18_stream_ivalid <= 0;
      end 
      case(__reduce_max_18_fsm)
        __reduce_max_18_fsm_init: begin
          if(__reduce_max_18_run_flag) begin
            __reduce_max_18_source_start <= 1;
          end 
          if(__reduce_max_18_run_flag) begin
            __reduce_max_18_fsm <= __reduce_max_18_fsm_1;
          end 
        end
        __reduce_max_18_fsm_1: begin
          if(__reduce_max_18_source_start && __reduce_max_18_stream_oready) begin
            __reduce_max_18_source_start <= 0;
            __reduce_max_18_source_busy <= 1;
          end 
          if(__reduce_max_18_source_start && __reduce_max_18_stream_oready) begin
            __reduce_max_18_fsm <= __reduce_max_18_fsm_2;
          end 
        end
        __reduce_max_18_fsm_2: begin
          if(__reduce_max_18_stream_oready) begin
            __reduce_max_18_fsm <= __reduce_max_18_fsm_3;
          end 
        end
        __reduce_max_18_fsm_3: begin
          if(__reduce_max_18_stream_oready && 1'd0) begin
            __reduce_max_18_source_busy <= 0;
          end 
          if(__reduce_max_18_stream_oready && 1'd0 && __reduce_max_18_run_flag) begin
            __reduce_max_18_source_start <= 1;
          end 
          if(__reduce_max_18_stream_oready && 1'd0) begin
            __reduce_max_18_fsm <= __reduce_max_18_fsm_init;
          end 
          if(__reduce_max_18_stream_oready && 1'd0 && __reduce_max_18_run_flag) begin
            __reduce_max_18_fsm <= __reduce_max_18_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_7_source_ram_renable <= 0;
      _stream_conv2d_4_source_7_source_fifo_deq <= 0;
      _stream_conv2d_4_source_7_idle <= 1;
      _stream_conv2d_4_source_9_source_ram_renable <= 0;
      _stream_conv2d_4_source_9_source_fifo_deq <= 0;
      _stream_conv2d_4_source_9_idle <= 1;
      _stream_conv2d_4_source_11_source_ram_renable <= 0;
      _stream_conv2d_4_source_11_source_fifo_deq <= 0;
      _stream_conv2d_4_source_11_idle <= 1;
      _stream_conv2d_4_source_13_source_ram_renable <= 0;
      _stream_conv2d_4_source_13_source_fifo_deq <= 0;
      _stream_conv2d_4_source_13_idle <= 1;
      _stream_conv2d_4_source_15_source_ram_renable <= 0;
      _stream_conv2d_4_source_15_source_fifo_deq <= 0;
      _stream_conv2d_4_source_15_idle <= 1;
      _stream_conv2d_4_source_20_source_ram_renable <= 0;
      _stream_conv2d_4_source_20_source_fifo_deq <= 0;
      _stream_conv2d_4_source_20_idle <= 1;
      _stream_conv2d_4_source_21_source_ram_renable <= 0;
      _stream_conv2d_4_source_21_source_fifo_deq <= 0;
      _stream_conv2d_4_source_21_idle <= 1;
      _stream_conv2d_4_source_22_source_ram_renable <= 0;
      _stream_conv2d_4_source_22_source_fifo_deq <= 0;
      _stream_conv2d_4_source_22_idle <= 1;
      _stream_conv2d_4_source_23_source_ram_renable <= 0;
      _stream_conv2d_4_source_23_source_fifo_deq <= 0;
      _stream_conv2d_4_source_23_idle <= 1;
      _stream_conv2d_4_source_24_source_ram_renable <= 0;
      _stream_conv2d_4_source_24_source_fifo_deq <= 0;
      _stream_conv2d_4_source_24_idle <= 1;
      _stream_conv2d_4_source_25_source_ram_renable <= 0;
      _stream_conv2d_4_source_25_source_fifo_deq <= 0;
      _stream_conv2d_4_source_25_idle <= 1;
      _stream_conv2d_4_source_26_source_ram_renable <= 0;
      _stream_conv2d_4_source_26_source_fifo_deq <= 0;
      _stream_conv2d_4_source_26_idle <= 1;
      _stream_conv2d_4_source_27_source_ram_renable <= 0;
      _stream_conv2d_4_source_27_source_fifo_deq <= 0;
      _stream_conv2d_4_source_27_idle <= 1;
      _stream_conv2d_4_source_28_source_ram_renable <= 0;
      _stream_conv2d_4_source_28_source_fifo_deq <= 0;
      _stream_conv2d_4_source_28_idle <= 1;
      _stream_conv2d_4_source_29_source_ram_renable <= 0;
      _stream_conv2d_4_source_29_source_fifo_deq <= 0;
      _stream_conv2d_4_source_29_idle <= 1;
      _stream_conv2d_4_source_30_source_ram_renable <= 0;
      _stream_conv2d_4_source_30_source_fifo_deq <= 0;
      _stream_conv2d_4_source_30_idle <= 1;
      _stream_conv2d_4_source_31_source_ram_renable <= 0;
      _stream_conv2d_4_source_31_source_fifo_deq <= 0;
      _stream_conv2d_4_source_31_idle <= 1;
      _stream_conv2d_4_source_32_source_ram_renable <= 0;
      _stream_conv2d_4_source_32_source_fifo_deq <= 0;
      _stream_conv2d_4_source_32_idle <= 1;
      _stream_conv2d_4_source_33_source_ram_renable <= 0;
      _stream_conv2d_4_source_33_source_fifo_deq <= 0;
      _stream_conv2d_4_source_33_idle <= 1;
      _stream_conv2d_4_source_34_source_ram_renable <= 0;
      _stream_conv2d_4_source_34_source_fifo_deq <= 0;
      _stream_conv2d_4_source_34_idle <= 1;
      _stream_conv2d_4_source_35_source_ram_renable <= 0;
      _stream_conv2d_4_source_35_source_fifo_deq <= 0;
      _stream_conv2d_4_source_35_idle <= 1;
      _stream_conv2d_4_source_36_source_ram_renable <= 0;
      _stream_conv2d_4_source_36_source_fifo_deq <= 0;
      _stream_conv2d_4_source_36_idle <= 1;
      _stream_conv2d_4_source_37_source_ram_renable <= 0;
      _stream_conv2d_4_source_37_source_fifo_deq <= 0;
      _stream_conv2d_4_source_37_idle <= 1;
      _stream_conv2d_4_sink_50_sink_wenable <= 0;
      _stream_conv2d_4_sink_50_sink_fifo_enq <= 0;
      _stream_conv2d_4_sink_51_sink_wenable <= 0;
      _stream_conv2d_4_sink_51_sink_fifo_enq <= 0;
      __stream_conv2d_4_stream_ivalid_1 <= 0;
      __stream_conv2d_4_stream_ivalid_2 <= 0;
      __stream_conv2d_4_stream_ivalid_3 <= 0;
      __stream_conv2d_4_stream_ivalid_4 <= 0;
      __stream_conv2d_4_stream_ivalid_5 <= 0;
      __stream_conv2d_4_stream_ivalid_6 <= 0;
      __stream_conv2d_4_stream_ivalid_7 <= 0;
      __stream_conv2d_4_stream_ivalid_8 <= 0;
      __stream_conv2d_4_stream_ivalid_9 <= 0;
      __stream_conv2d_4_stream_ivalid_10 <= 0;
      __stream_conv2d_4_stream_ivalid_11 <= 0;
      __stream_conv2d_4_stream_ivalid_12 <= 0;
      __stream_conv2d_4_stream_ivalid_13 <= 0;
      __stream_conv2d_4_stream_ivalid_14 <= 0;
      __stream_conv2d_4_stream_ivalid_15 <= 0;
      __stream_conv2d_4_stream_ivalid_16 <= 0;
      __stream_conv2d_4_stream_ivalid_17 <= 0;
      __stream_conv2d_4_stream_ivalid_18 <= 0;
      __stream_conv2d_4_stream_ivalid_19 <= 0;
      __stream_conv2d_4_stream_ivalid_20 <= 0;
      __stream_conv2d_4_stream_ivalid_21 <= 0;
      __stream_conv2d_4_stream_ivalid_22 <= 0;
      __stream_conv2d_4_stream_ivalid_23 <= 0;
      __stream_conv2d_4_stream_ivalid_24 <= 0;
      __stream_conv2d_4_stream_ivalid_25 <= 0;
      __stream_conv2d_4_stream_ivalid_26 <= 0;
      __stream_conv2d_4_stream_ivalid_27 <= 0;
      __stream_conv2d_4_stream_ivalid_28 <= 0;
      __stream_conv2d_4_stream_ivalid_29 <= 0;
      __stream_conv2d_4_stream_ivalid_30 <= 0;
      __stream_conv2d_4_stream_ivalid_31 <= 0;
      _eq_data_402 <= 0;
      _eq_data_406 <= 0;
      _eq_data_409 <= 0;
      _eq_data_412 <= 0;
      _eq_data_416 <= 0;
      _eq_data_419 <= 0;
      _eq_data_422 <= 0;
      _eq_data_426 <= 0;
      _eq_data_429 <= 0;
      _eq_data_432 <= 0;
      _eq_data_436 <= 0;
      _eq_data_439 <= 0;
      _eq_data_442 <= 0;
      _eq_data_446 <= 0;
      _eq_data_449 <= 0;
      _eq_data_452 <= 0;
      _eq_data_456 <= 0;
      _eq_data_459 <= 0;
      _eq_data_462 <= 0;
      _eq_data_466 <= 0;
      _eq_data_469 <= 0;
      _eq_data_472 <= 0;
      _eq_data_476 <= 0;
      _eq_data_479 <= 0;
      _eq_data_482 <= 0;
      _eq_data_486 <= 0;
      _eq_data_489 <= 0;
      _eq_data_492 <= 0;
      _eq_data_496 <= 0;
      _eq_data_499 <= 0;
      _eq_data_502 <= 0;
      _eq_data_506 <= 0;
      _eq_data_509 <= 0;
      _eq_data_512 <= 0;
      _eq_data_516 <= 0;
      _eq_data_519 <= 0;
      _eq_data_522 <= 0;
      _eq_data_526 <= 0;
      _eq_data_529 <= 0;
      _eq_data_532 <= 0;
      _eq_data_536 <= 0;
      _eq_data_539 <= 0;
      _eq_data_542 <= 0;
      _eq_data_546 <= 0;
      _eq_data_549 <= 0;
      _eq_data_552 <= 0;
      _eq_data_556 <= 0;
      _eq_data_559 <= 0;
      _eq_data_562 <= 0;
      _eq_data_566 <= 0;
      _eq_data_569 <= 0;
      _eq_data_572 <= 0;
      _eq_data_576 <= 0;
      _eq_data_579 <= 0;
      _plus_data_734 <= 0;
      _plus_data_753 <= 0;
      _plus_data_772 <= 0;
      _plus_data_791 <= 0;
      _plus_data_810 <= 0;
      _plus_data_829 <= 0;
      _plus_data_848 <= 0;
      _plus_data_867 <= 0;
      _plus_data_886 <= 0;
      _plus_data_902 <= 0;
      _plus_data_921 <= 0;
      __delay_data_1254__variable_395 <= 0;
      __delay_data_1255__variable_394 <= 0;
      __delay_data_1256__variable_393 <= 0;
      __delay_data_1257__variable_398 <= 0;
      __delay_data_1258__variable_397 <= 0;
      __delay_data_1259__variable_396 <= 0;
      __delay_data_1260__variable_401 <= 0;
      __delay_data_1261__variable_400 <= 0;
      __delay_data_1262__variable_399 <= 0;
      __delay_data_1263_pointer_681 <= 0;
      __delay_data_1264_reinterpretcast_672 <= 0;
      __delay_data_1265_pointer_683 <= 0;
      __delay_data_1266_reinterpretcast_673 <= 0;
      __delay_data_1267_pointer_685 <= 0;
      __delay_data_1268_reinterpretcast_674 <= 0;
      __delay_data_1269_pointer_687 <= 0;
      __delay_data_1270_reinterpretcast_675 <= 0;
      __delay_data_1271_pointer_689 <= 0;
      __delay_data_1272_reinterpretcast_676 <= 0;
      __delay_data_1273_pointer_691 <= 0;
      __delay_data_1274_reinterpretcast_677 <= 0;
      __delay_data_1275_pointer_693 <= 0;
      __delay_data_1276_reinterpretcast_678 <= 0;
      __delay_data_1277_pointer_695 <= 0;
      __delay_data_1278_reinterpretcast_679 <= 0;
      __delay_data_1279_pointer_697 <= 0;
      __delay_data_1280_reinterpretcast_680 <= 0;
      __delay_data_1281__variable_344 <= 0;
      __delay_data_1306__variable_339 <= 0;
      __delay_data_1319_cond_360 <= 0;
      __delay_data_1338_cond_367 <= 0;
      __delay_data_1282__delay_1281__variable_344 <= 0;
      __delay_data_1294_plus_902 <= 0;
      __delay_data_1307__delay_1306__variable_339 <= 0;
      __delay_data_1320__delay_1319_cond_360 <= 0;
      __delay_data_1339__delay_1338_cond_367 <= 0;
      __delay_data_1358_plus_921 <= 0;
      __delay_data_1283__delay_1282__delay_1281__variable_344 <= 0;
      __delay_data_1295__delay_1294_plus_902 <= 0;
      __delay_data_1308__delay_1307__delay_1306__variable_339 <= 0;
      __delay_data_1321__delay_1320__delay_1319_cond_360 <= 0;
      __delay_data_1340__delay_1339__delay_1338_cond_367 <= 0;
      __delay_data_1359__delay_1358_plus_921 <= 0;
      __delay_data_1284__delay_1283__delay_1282____variable_344 <= 0;
      __delay_data_1296__delay_1295__delay_1294_plus_902 <= 0;
      __delay_data_1309__delay_1308__delay_1307____variable_339 <= 0;
      __delay_data_1322__delay_1321__delay_1320__delay_1319_cond_360 <= 0;
      __delay_data_1341__delay_1340__delay_1339__delay_1338_cond_367 <= 0;
      __delay_data_1360__delay_1359__delay_1358_plus_921 <= 0;
      __delay_data_1285__delay_1284__delay_1283____variable_344 <= 0;
      __delay_data_1297__delay_1296__delay_1295__delay_1294_plus_902 <= 0;
      __delay_data_1310__delay_1309__delay_1308____variable_339 <= 0;
      __delay_data_1323__delay_1322__delay_1321__delay_1320___cond_360 <= 0;
      __delay_data_1342__delay_1341__delay_1340__delay_1339___cond_367 <= 0;
      __delay_data_1361__delay_1360__delay_1359__delay_1358_plus_921 <= 0;
      __delay_data_1286__delay_1285__delay_1284____variable_344 <= 0;
      __delay_data_1298__delay_1297__delay_1296__delay_1295___plus_902 <= 0;
      __delay_data_1311__delay_1310__delay_1309____variable_339 <= 0;
      __delay_data_1324__delay_1323__delay_1322__delay_1321___cond_360 <= 0;
      __delay_data_1343__delay_1342__delay_1341__delay_1340___cond_367 <= 0;
      __delay_data_1362__delay_1361__delay_1360__delay_1359___plus_921 <= 0;
      __delay_data_1287__delay_1286__delay_1285____variable_344 <= 0;
      __delay_data_1299__delay_1298__delay_1297__delay_1296___plus_902 <= 0;
      __delay_data_1312__delay_1311__delay_1310____variable_339 <= 0;
      __delay_data_1325__delay_1324__delay_1323__delay_1322___cond_360 <= 0;
      __delay_data_1344__delay_1343__delay_1342__delay_1341___cond_367 <= 0;
      __delay_data_1363__delay_1362__delay_1361__delay_1360___plus_921 <= 0;
      __delay_data_1288__delay_1287__delay_1286____variable_344 <= 0;
      __delay_data_1300__delay_1299__delay_1298__delay_1297___plus_902 <= 0;
      __delay_data_1313__delay_1312__delay_1311____variable_339 <= 0;
      __delay_data_1326__delay_1325__delay_1324__delay_1323___cond_360 <= 0;
      __delay_data_1345__delay_1344__delay_1343__delay_1342___cond_367 <= 0;
      __delay_data_1364__delay_1363__delay_1362__delay_1361___plus_921 <= 0;
      __delay_data_1289__delay_1288__delay_1287____variable_344 <= 0;
      __delay_data_1301__delay_1300__delay_1299__delay_1298___plus_902 <= 0;
      __delay_data_1314__delay_1313__delay_1312____variable_339 <= 0;
      __delay_data_1327__delay_1326__delay_1325__delay_1324___cond_360 <= 0;
      __delay_data_1346__delay_1345__delay_1344__delay_1343___cond_367 <= 0;
      __delay_data_1365__delay_1364__delay_1363__delay_1362___plus_921 <= 0;
      __delay_data_1290__delay_1289__delay_1288____variable_344 <= 0;
      __delay_data_1302__delay_1301__delay_1300__delay_1299___plus_902 <= 0;
      __delay_data_1315__delay_1314__delay_1313____variable_339 <= 0;
      __delay_data_1328__delay_1327__delay_1326__delay_1325___cond_360 <= 0;
      __delay_data_1347__delay_1346__delay_1345__delay_1344___cond_367 <= 0;
      __delay_data_1366__delay_1365__delay_1364__delay_1363___plus_921 <= 0;
      __delay_data_1291__delay_1290__delay_1289____variable_344 <= 0;
      __delay_data_1303__delay_1302__delay_1301__delay_1300___plus_902 <= 0;
      __delay_data_1316__delay_1315__delay_1314____variable_339 <= 0;
      __delay_data_1329__delay_1328__delay_1327__delay_1326___cond_360 <= 0;
      __delay_data_1348__delay_1347__delay_1346__delay_1345___cond_367 <= 0;
      __delay_data_1367__delay_1366__delay_1365__delay_1364___plus_921 <= 0;
      __delay_data_1292__delay_1291__delay_1290____variable_344 <= 0;
      __delay_data_1304__delay_1303__delay_1302__delay_1301___plus_902 <= 0;
      __delay_data_1317__delay_1316__delay_1315____variable_339 <= 0;
      __delay_data_1330__delay_1329__delay_1328__delay_1327___cond_360 <= 0;
      __delay_data_1349__delay_1348__delay_1347__delay_1346___cond_367 <= 0;
      __delay_data_1368__delay_1367__delay_1366__delay_1365___plus_921 <= 0;
      __delay_data_1293__delay_1292__delay_1291____variable_344 <= 0;
      __delay_data_1305__delay_1304__delay_1303__delay_1302___plus_902 <= 0;
      __delay_data_1318__delay_1317__delay_1316____variable_339 <= 0;
      __delay_data_1331__delay_1330__delay_1329__delay_1328___cond_360 <= 0;
      __delay_data_1350__delay_1349__delay_1348__delay_1347___cond_367 <= 0;
      __delay_data_1369__delay_1368__delay_1367__delay_1366___plus_921 <= 0;
      __delay_data_1332__delay_1331__delay_1330__delay_1329___cond_360 <= 0;
      __delay_data_1351__delay_1350__delay_1349__delay_1348___cond_367 <= 0;
      __delay_data_1370__delay_1369__delay_1368__delay_1367___plus_921 <= 0;
      __delay_data_1333__delay_1332__delay_1331__delay_1330___cond_360 <= 0;
      __delay_data_1352__delay_1351__delay_1350__delay_1349___cond_367 <= 0;
      __delay_data_1371__delay_1370__delay_1369__delay_1368___plus_921 <= 0;
      __delay_data_1334__delay_1333__delay_1332__delay_1331___cond_360 <= 0;
      __delay_data_1353__delay_1352__delay_1351__delay_1350___cond_367 <= 0;
      __delay_data_1372__delay_1371__delay_1370__delay_1369___plus_921 <= 0;
      __delay_data_1335__delay_1334__delay_1333__delay_1332___cond_360 <= 0;
      __delay_data_1354__delay_1353__delay_1352__delay_1351___cond_367 <= 0;
      __delay_data_1373__delay_1372__delay_1371__delay_1370___plus_921 <= 0;
      __delay_data_1336__delay_1335__delay_1334__delay_1333___cond_360 <= 0;
      __delay_data_1355__delay_1354__delay_1353__delay_1352___cond_367 <= 0;
      __delay_data_1374__delay_1373__delay_1372__delay_1371___plus_921 <= 0;
      __delay_data_1337__delay_1336__delay_1335__delay_1334___cond_360 <= 0;
      __delay_data_1356__delay_1355__delay_1354__delay_1353___cond_367 <= 0;
      __delay_data_1375__delay_1374__delay_1373__delay_1372___plus_921 <= 0;
      _plus_data_905 <= 0;
      __delay_data_1357__delay_1356__delay_1355__delay_1354___cond_367 <= 0;
      __delay_data_1376__delay_1375__delay_1374__delay_1373___plus_921 <= 0;
      __delay_data_1378__substreamoutput_904 <= 0;
      __delay_data_1379__delay_1378__substreamoutput_904 <= 0;
      __delay_data_1380__delay_1379__delay_1378__substreamoutput_904 <= 0;
      __delay_data_1381__delay_1380__delay_1379____substreamoutput_904 <= 0;
      __delay_data_1382__delay_1381__delay_1380____substreamoutput_904 <= 0;
      __delay_data_1383__delay_1382__delay_1381____substreamoutput_904 <= 0;
      __delay_data_1384__delay_1383__delay_1382____substreamoutput_904 <= 0;
      __delay_data_1385__delay_1384__delay_1383____substreamoutput_904 <= 0;
      __delay_data_1386__delay_1385__delay_1384____substreamoutput_904 <= 0;
      __delay_data_1387__delay_1386__delay_1385____substreamoutput_904 <= 0;
      _greaterthan_data_924 <= 0;
      __delay_data_1377__substreamoutput_922 <= 0;
      __delay_data_1388__delay_1387__delay_1386____substreamoutput_904 <= 0;
      _cond_data_926 <= 0;
      __delay_data_1389__delay_1388__delay_1387____substreamoutput_904 <= 0;
      _stream_conv2d_4_parameter_0_next_parameter_data <= 0;
      __variable_wdata_339 <= 0;
      _stream_conv2d_4_parameter_1_next_parameter_data <= 0;
      __variable_wdata_340 <= 0;
      _stream_conv2d_4_parameter_2_next_parameter_data <= 0;
      __variable_wdata_341 <= 0;
      _stream_conv2d_4_parameter_3_next_parameter_data <= 0;
      __variable_wdata_342 <= 0;
      _stream_conv2d_4_parameter_4_next_parameter_data <= 0;
      __variable_wdata_343 <= 0;
      _stream_conv2d_4_parameter_6_next_parameter_data <= 0;
      __variable_wdata_354 <= 0;
      _stream_conv2d_4_source_7_source_mode <= 5'b0;
      _stream_conv2d_4_source_7_source_offset <= 0;
      _source_stream_conv2d_4_source_7_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_3 <= 0;
      _stream_conv2d_4_source_7_source_sel <= 0;
      _stream_conv2d_4_source_7_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_7_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_7_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_buf_3 <= 0;
      __variable_wdata_355 <= 0;
      _stream_conv2d_4_source_7_source_ram_raddr <= 0;
      _stream_conv2d_4_parameter_8_next_parameter_data <= 0;
      __variable_wdata_361 <= 0;
      _stream_conv2d_4_source_9_source_mode <= 5'b0;
      _stream_conv2d_4_source_9_source_offset <= 0;
      _source_stream_conv2d_4_source_9_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_3 <= 0;
      _stream_conv2d_4_source_9_source_sel <= 0;
      _stream_conv2d_4_source_9_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_9_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_9_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_buf_3 <= 0;
      __variable_wdata_362 <= 0;
      _stream_conv2d_4_source_9_source_ram_raddr <= 0;
      _stream_conv2d_4_parameter_10_next_parameter_data <= 0;
      __variable_wdata_368 <= 0;
      _stream_conv2d_4_source_11_source_mode <= 5'b0;
      _stream_conv2d_4_source_11_source_empty_data <= 0;
      __variable_wdata_369 <= 0;
      _stream_conv2d_4_parameter_12_next_parameter_data <= 0;
      __variable_wdata_375 <= 0;
      _stream_conv2d_4_source_13_source_mode <= 5'b0;
      _stream_conv2d_4_source_13_source_empty_data <= 0;
      __variable_wdata_376 <= 0;
      _stream_conv2d_4_parameter_14_next_parameter_data <= 0;
      __variable_wdata_382 <= 0;
      _stream_conv2d_4_source_15_source_mode <= 5'b0;
      _stream_conv2d_4_source_15_source_empty_data <= 0;
      __variable_wdata_383 <= 0;
      _stream_conv2d_4_parameter_16_next_parameter_data <= 0;
      __variable_wdata_389 <= 0;
      _stream_conv2d_4_parameter_17_next_parameter_data <= 0;
      __variable_wdata_390 <= 0;
      _stream_conv2d_4_parameter_18_next_parameter_data <= 0;
      __variable_wdata_391 <= 0;
      _stream_conv2d_4_parameter_19_next_parameter_data <= 0;
      __variable_wdata_392 <= 0;
      _stream_conv2d_4_source_20_source_mode <= 5'b0;
      _stream_conv2d_4_source_20_source_offset <= 0;
      _source_stream_conv2d_4_source_20_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_3 <= 0;
      _stream_conv2d_4_source_20_source_sel <= 0;
      _stream_conv2d_4_source_20_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_20_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_20_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_buf_3 <= 0;
      __variable_wdata_393 <= 0;
      _stream_conv2d_4_source_20_source_ram_raddr <= 0;
      _stream_conv2d_4_source_21_source_mode <= 5'b0;
      _stream_conv2d_4_source_21_source_offset <= 0;
      _source_stream_conv2d_4_source_21_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_3 <= 0;
      _stream_conv2d_4_source_21_source_sel <= 0;
      _stream_conv2d_4_source_21_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_21_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_21_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_buf_3 <= 0;
      __variable_wdata_394 <= 0;
      _stream_conv2d_4_source_21_source_ram_raddr <= 0;
      _stream_conv2d_4_source_22_source_mode <= 5'b0;
      _stream_conv2d_4_source_22_source_offset <= 0;
      _source_stream_conv2d_4_source_22_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_3 <= 0;
      _stream_conv2d_4_source_22_source_sel <= 0;
      _stream_conv2d_4_source_22_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_22_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_22_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_buf_3 <= 0;
      __variable_wdata_395 <= 0;
      _stream_conv2d_4_source_22_source_ram_raddr <= 0;
      _stream_conv2d_4_source_23_source_mode <= 5'b0;
      _stream_conv2d_4_source_23_source_offset <= 0;
      _source_stream_conv2d_4_source_23_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_3 <= 0;
      _stream_conv2d_4_source_23_source_sel <= 0;
      _stream_conv2d_4_source_23_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_23_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_23_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_buf_3 <= 0;
      __variable_wdata_396 <= 0;
      _stream_conv2d_4_source_23_source_ram_raddr <= 0;
      _stream_conv2d_4_source_24_source_mode <= 5'b0;
      _stream_conv2d_4_source_24_source_offset <= 0;
      _source_stream_conv2d_4_source_24_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_3 <= 0;
      _stream_conv2d_4_source_24_source_sel <= 0;
      _stream_conv2d_4_source_24_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_24_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_24_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_buf_3 <= 0;
      __variable_wdata_397 <= 0;
      _stream_conv2d_4_source_24_source_ram_raddr <= 0;
      _stream_conv2d_4_source_25_source_mode <= 5'b0;
      _stream_conv2d_4_source_25_source_offset <= 0;
      _source_stream_conv2d_4_source_25_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_3 <= 0;
      _stream_conv2d_4_source_25_source_sel <= 0;
      _stream_conv2d_4_source_25_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_25_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_25_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_buf_3 <= 0;
      __variable_wdata_398 <= 0;
      _stream_conv2d_4_source_25_source_ram_raddr <= 0;
      _stream_conv2d_4_source_26_source_mode <= 5'b0;
      _stream_conv2d_4_source_26_source_offset <= 0;
      _source_stream_conv2d_4_source_26_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_3 <= 0;
      _stream_conv2d_4_source_26_source_sel <= 0;
      _stream_conv2d_4_source_26_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_26_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_26_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_buf_3 <= 0;
      __variable_wdata_399 <= 0;
      _stream_conv2d_4_source_26_source_ram_raddr <= 0;
      _stream_conv2d_4_source_27_source_mode <= 5'b0;
      _stream_conv2d_4_source_27_source_offset <= 0;
      _source_stream_conv2d_4_source_27_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_3 <= 0;
      _stream_conv2d_4_source_27_source_sel <= 0;
      _stream_conv2d_4_source_27_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_27_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_27_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_buf_3 <= 0;
      __variable_wdata_400 <= 0;
      _stream_conv2d_4_source_27_source_ram_raddr <= 0;
      _stream_conv2d_4_source_28_source_mode <= 5'b0;
      _stream_conv2d_4_source_28_source_offset <= 0;
      _source_stream_conv2d_4_source_28_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_3 <= 0;
      _stream_conv2d_4_source_28_source_sel <= 0;
      _stream_conv2d_4_source_28_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_28_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_28_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_buf_3 <= 0;
      __variable_wdata_401 <= 0;
      _stream_conv2d_4_source_28_source_ram_raddr <= 0;
      _stream_conv2d_4_source_29_source_mode <= 5'b0;
      _stream_conv2d_4_source_29_source_offset <= 0;
      _source_stream_conv2d_4_source_29_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_3 <= 0;
      _stream_conv2d_4_source_29_source_sel <= 0;
      _stream_conv2d_4_source_29_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_29_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_29_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_buf_3 <= 0;
      __variable_wdata_627 <= 0;
      _stream_conv2d_4_source_29_source_ram_raddr <= 0;
      _stream_conv2d_4_source_30_source_mode <= 5'b0;
      _stream_conv2d_4_source_30_source_offset <= 0;
      _source_stream_conv2d_4_source_30_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_3 <= 0;
      _stream_conv2d_4_source_30_source_sel <= 0;
      _stream_conv2d_4_source_30_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_30_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_30_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_buf_3 <= 0;
      __variable_wdata_628 <= 0;
      _stream_conv2d_4_source_30_source_ram_raddr <= 0;
      _stream_conv2d_4_source_31_source_mode <= 5'b0;
      _stream_conv2d_4_source_31_source_offset <= 0;
      _source_stream_conv2d_4_source_31_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_3 <= 0;
      _stream_conv2d_4_source_31_source_sel <= 0;
      _stream_conv2d_4_source_31_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_31_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_31_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_buf_3 <= 0;
      __variable_wdata_629 <= 0;
      _stream_conv2d_4_source_31_source_ram_raddr <= 0;
      _stream_conv2d_4_source_32_source_mode <= 5'b0;
      _stream_conv2d_4_source_32_source_offset <= 0;
      _source_stream_conv2d_4_source_32_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_3 <= 0;
      _stream_conv2d_4_source_32_source_sel <= 0;
      _stream_conv2d_4_source_32_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_32_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_32_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_buf_3 <= 0;
      __variable_wdata_630 <= 0;
      _stream_conv2d_4_source_32_source_ram_raddr <= 0;
      _stream_conv2d_4_source_33_source_mode <= 5'b0;
      _stream_conv2d_4_source_33_source_offset <= 0;
      _source_stream_conv2d_4_source_33_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_3 <= 0;
      _stream_conv2d_4_source_33_source_sel <= 0;
      _stream_conv2d_4_source_33_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_33_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_33_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_buf_3 <= 0;
      __variable_wdata_631 <= 0;
      _stream_conv2d_4_source_33_source_ram_raddr <= 0;
      _stream_conv2d_4_source_34_source_mode <= 5'b0;
      _stream_conv2d_4_source_34_source_offset <= 0;
      _source_stream_conv2d_4_source_34_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_3 <= 0;
      _stream_conv2d_4_source_34_source_sel <= 0;
      _stream_conv2d_4_source_34_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_34_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_34_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_buf_3 <= 0;
      __variable_wdata_632 <= 0;
      _stream_conv2d_4_source_34_source_ram_raddr <= 0;
      _stream_conv2d_4_source_35_source_mode <= 5'b0;
      _stream_conv2d_4_source_35_source_offset <= 0;
      _source_stream_conv2d_4_source_35_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_3 <= 0;
      _stream_conv2d_4_source_35_source_sel <= 0;
      _stream_conv2d_4_source_35_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_35_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_35_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_buf_3 <= 0;
      __variable_wdata_633 <= 0;
      _stream_conv2d_4_source_35_source_ram_raddr <= 0;
      _stream_conv2d_4_source_36_source_mode <= 5'b0;
      _stream_conv2d_4_source_36_source_offset <= 0;
      _source_stream_conv2d_4_source_36_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_3 <= 0;
      _stream_conv2d_4_source_36_source_sel <= 0;
      _stream_conv2d_4_source_36_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_36_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_36_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_buf_3 <= 0;
      __variable_wdata_634 <= 0;
      _stream_conv2d_4_source_36_source_ram_raddr <= 0;
      _stream_conv2d_4_source_37_source_mode <= 5'b0;
      _stream_conv2d_4_source_37_source_offset <= 0;
      _source_stream_conv2d_4_source_37_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_3 <= 0;
      _stream_conv2d_4_source_37_source_sel <= 0;
      _stream_conv2d_4_source_37_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_37_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_37_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_buf_3 <= 0;
      __variable_wdata_635 <= 0;
      _stream_conv2d_4_source_37_source_ram_raddr <= 0;
      _tmp_526 <= 0;
      _tmp_527 <= 0;
      _tmp_528 <= 0;
      _tmp_529 <= 0;
      _tmp_530 <= 0;
      _tmp_531 <= 0;
      _tmp_532 <= 0;
      _tmp_533 <= 0;
      _tmp_534 <= 0;
      _tmp_535 <= 0;
      _tmp_536 <= 0;
      _tmp_537 <= 0;
      _tmp_538 <= 0;
      _tmp_539 <= 0;
      _tmp_540 <= 0;
      _tmp_541 <= 0;
      _tmp_542 <= 0;
      _tmp_543 <= 0;
      _tmp_544 <= 0;
      _tmp_545 <= 0;
      _tmp_546 <= 0;
      _tmp_547 <= 0;
      _tmp_548 <= 0;
      _tmp_549 <= 0;
      _tmp_550 <= 0;
      _tmp_551 <= 0;
      _tmp_552 <= 0;
      _tmp_553 <= 0;
      _tmp_554 <= 0;
      _tmp_555 <= 0;
      _tmp_556 <= 0;
      _tmp_557 <= 0;
      _tmp_558 <= 0;
      _tmp_561 <= 0;
      _tmp_562 <= 0;
      _tmp_563 <= 0;
      _tmp_564 <= 0;
      _tmp_565 <= 0;
      _tmp_566 <= 0;
      _tmp_567 <= 0;
      _tmp_568 <= 0;
      _tmp_569 <= 0;
      _tmp_570 <= 0;
      _tmp_571 <= 0;
      _tmp_572 <= 0;
      _tmp_573 <= 0;
      _tmp_574 <= 0;
      _tmp_575 <= 0;
      _tmp_576 <= 0;
      _tmp_577 <= 0;
      _tmp_578 <= 0;
      _tmp_579 <= 0;
      _tmp_580 <= 0;
      _tmp_581 <= 0;
      _tmp_582 <= 0;
      _tmp_583 <= 0;
      _tmp_584 <= 0;
      _tmp_585 <= 0;
      _tmp_586 <= 0;
      _tmp_587 <= 0;
      _tmp_588 <= 0;
      _tmp_589 <= 0;
      _tmp_590 <= 0;
      _tmp_591 <= 0;
      _tmp_592 <= 0;
      _tmp_593 <= 0;
      _tmp_594 <= 0;
      _tmp_595 <= 0;
      _tmp_596 <= 0;
      _tmp_597 <= 0;
      _tmp_598 <= 0;
      _tmp_599 <= 0;
      _tmp_600 <= 0;
      _tmp_601 <= 0;
      _tmp_602 <= 0;
      _tmp_603 <= 0;
      _tmp_604 <= 0;
      _tmp_605 <= 0;
      _tmp_606 <= 0;
      _tmp_607 <= 0;
      _tmp_608 <= 0;
      _tmp_609 <= 0;
      _tmp_610 <= 0;
      _tmp_611 <= 0;
      _tmp_612 <= 0;
      _tmp_613 <= 0;
      _tmp_614 <= 0;
      _tmp_615 <= 0;
      _tmp_616 <= 0;
      _tmp_617 <= 0;
      _tmp_618 <= 0;
      _tmp_619 <= 0;
      _tmp_620 <= 0;
      _tmp_621 <= 0;
      _tmp_622 <= 0;
      _tmp_623 <= 0;
      _tmp_624 <= 0;
      _tmp_625 <= 0;
      _tmp_626 <= 0;
      _stream_conv2d_4_sink_50_sink_mode <= 5'b0;
      _stream_conv2d_4_sink_50_sink_offset <= 0;
      _stream_conv2d_4_sink_50_sink_size <= 0;
      _stream_conv2d_4_sink_50_sink_stride <= 0;
      _stream_conv2d_4_sink_50_sink_sel <= 0;
      _stream_conv2d_4_sink_50_sink_offset_buf <= 0;
      _stream_conv2d_4_sink_50_sink_size_buf <= 0;
      _stream_conv2d_4_sink_50_sink_stride_buf <= 0;
      _stream_conv2d_4_sink_50_sink_waddr <= 0;
      _stream_conv2d_4_sink_50_sink_count <= 0;
      _stream_conv2d_4_sink_50_sink_wdata <= 0;
      _tmp_1017 <= 0;
      _tmp_1018 <= 0;
      _tmp_1019 <= 0;
      _tmp_1020 <= 0;
      _tmp_1021 <= 0;
      _tmp_1022 <= 0;
      __variable_wdata_344 <= 0;
      _tmp_1023 <= 0;
      _tmp_1024 <= 0;
      _tmp_1025 <= 0;
      _tmp_1026 <= 0;
      _tmp_1029 <= 0;
      _tmp_1032 <= 0;
      _tmp_1033 <= 0;
      _tmp_1034 <= 0;
      _tmp_1035 <= 0;
      _tmp_1036 <= 0;
      _tmp_1037 <= 0;
      _tmp_1038 <= 0;
      _tmp_1039 <= 0;
      _tmp_1040 <= 0;
      _tmp_1041 <= 0;
      _tmp_1042 <= 0;
      _tmp_1043 <= 0;
      _tmp_1044 <= 0;
      _tmp_1045 <= 0;
      _tmp_1046 <= 0;
      _tmp_1047 <= 0;
      _tmp_1048 <= 0;
      _tmp_1049 <= 0;
      _tmp_1050 <= 0;
      _tmp_1051 <= 0;
      _tmp_1052 <= 0;
      _tmp_1053 <= 0;
      _tmp_1054 <= 0;
      _tmp_1055 <= 0;
      _tmp_1056 <= 0;
      _tmp_1057 <= 0;
      _tmp_1058 <= 0;
      _tmp_1059 <= 0;
      _tmp_1060 <= 0;
      _tmp_1061 <= 0;
      _tmp_1062 <= 0;
      _tmp_1063 <= 0;
      _tmp_1064 <= 0;
      _tmp_1065 <= 0;
      _tmp_1066 <= 0;
      _tmp_1067 <= 0;
      _tmp_1068 <= 0;
      _tmp_1069 <= 0;
      _tmp_1070 <= 0;
      _tmp_1071 <= 0;
      _tmp_1072 <= 0;
      _tmp_1073 <= 0;
      _tmp_1074 <= 0;
      _tmp_1075 <= 0;
      _tmp_1076 <= 0;
      _tmp_1077 <= 0;
      _tmp_1078 <= 0;
      _tmp_1079 <= 0;
      _tmp_1080 <= 0;
      _tmp_1081 <= 0;
      _tmp_1082 <= 0;
      _tmp_1083 <= 0;
      _tmp_1084 <= 0;
      _tmp_1085 <= 0;
      _tmp_1086 <= 0;
      _tmp_1087 <= 0;
      _tmp_1088 <= 0;
      _tmp_1089 <= 0;
      _tmp_1090 <= 0;
      _tmp_1091 <= 0;
      _tmp_1092 <= 0;
      _tmp_1093 <= 0;
      _tmp_1094 <= 0;
      _tmp_1095 <= 0;
      _tmp_1096 <= 0;
      _tmp_1097 <= 0;
      _tmp_1098 <= 0;
      _tmp_1099 <= 0;
      _tmp_1100 <= 0;
      _tmp_1101 <= 0;
      _tmp_1102 <= 0;
      _tmp_1103 <= 0;
      _tmp_1104 <= 0;
      _tmp_1105 <= 0;
      _tmp_1106 <= 0;
      _tmp_1107 <= 0;
      _tmp_1108 <= 0;
      _tmp_1109 <= 0;
      _tmp_1110 <= 0;
      _tmp_1111 <= 0;
      _tmp_1112 <= 0;
      _tmp_1113 <= 0;
      _tmp_1114 <= 0;
      _tmp_1115 <= 0;
      _tmp_1116 <= 0;
      _tmp_1117 <= 0;
      _tmp_1118 <= 0;
      _tmp_1119 <= 0;
      _tmp_1120 <= 0;
      _tmp_1121 <= 0;
      _tmp_1122 <= 0;
      _tmp_1123 <= 0;
      _tmp_1124 <= 0;
      _tmp_1125 <= 0;
      _tmp_1126 <= 0;
      _tmp_1127 <= 0;
      _tmp_1128 <= 0;
      _tmp_1129 <= 0;
      _tmp_1130 <= 0;
      _tmp_1131 <= 0;
      _tmp_1132 <= 0;
      _stream_conv2d_4_busy_reg <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_source_ram_renable <= 0;
        _stream_conv2d_4_source_7_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_7_idle <= _stream_conv2d_4_source_7_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_source_ram_renable <= 0;
        _stream_conv2d_4_source_9_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_9_idle <= _stream_conv2d_4_source_9_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_11_source_ram_renable <= 0;
        _stream_conv2d_4_source_11_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_11_idle <= _stream_conv2d_4_source_11_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_13_source_ram_renable <= 0;
        _stream_conv2d_4_source_13_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_13_idle <= _stream_conv2d_4_source_13_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_15_source_ram_renable <= 0;
        _stream_conv2d_4_source_15_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_15_idle <= _stream_conv2d_4_source_15_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_source_ram_renable <= 0;
        _stream_conv2d_4_source_20_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_20_idle <= _stream_conv2d_4_source_20_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_source_ram_renable <= 0;
        _stream_conv2d_4_source_21_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_21_idle <= _stream_conv2d_4_source_21_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_source_ram_renable <= 0;
        _stream_conv2d_4_source_22_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_22_idle <= _stream_conv2d_4_source_22_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_source_ram_renable <= 0;
        _stream_conv2d_4_source_23_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_23_idle <= _stream_conv2d_4_source_23_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_source_ram_renable <= 0;
        _stream_conv2d_4_source_24_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_24_idle <= _stream_conv2d_4_source_24_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_source_ram_renable <= 0;
        _stream_conv2d_4_source_25_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_25_idle <= _stream_conv2d_4_source_25_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_source_ram_renable <= 0;
        _stream_conv2d_4_source_26_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_26_idle <= _stream_conv2d_4_source_26_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_source_ram_renable <= 0;
        _stream_conv2d_4_source_27_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_27_idle <= _stream_conv2d_4_source_27_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_source_ram_renable <= 0;
        _stream_conv2d_4_source_28_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_28_idle <= _stream_conv2d_4_source_28_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_source_ram_renable <= 0;
        _stream_conv2d_4_source_29_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_29_idle <= _stream_conv2d_4_source_29_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_source_ram_renable <= 0;
        _stream_conv2d_4_source_30_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_30_idle <= _stream_conv2d_4_source_30_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_source_ram_renable <= 0;
        _stream_conv2d_4_source_31_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_31_idle <= _stream_conv2d_4_source_31_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_source_ram_renable <= 0;
        _stream_conv2d_4_source_32_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_32_idle <= _stream_conv2d_4_source_32_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_source_ram_renable <= 0;
        _stream_conv2d_4_source_33_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_33_idle <= _stream_conv2d_4_source_33_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_source_ram_renable <= 0;
        _stream_conv2d_4_source_34_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_34_idle <= _stream_conv2d_4_source_34_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_source_ram_renable <= 0;
        _stream_conv2d_4_source_35_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_35_idle <= _stream_conv2d_4_source_35_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_source_ram_renable <= 0;
        _stream_conv2d_4_source_36_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_36_idle <= _stream_conv2d_4_source_36_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_source_ram_renable <= 0;
        _stream_conv2d_4_source_37_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_37_idle <= _stream_conv2d_4_source_37_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_50_sink_wenable <= 0;
        _stream_conv2d_4_sink_50_sink_fifo_enq <= 0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_51_sink_wenable <= 0;
        _stream_conv2d_4_sink_51_sink_fifo_enq <= 0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_1 <= _stream_conv2d_4_stream_ivalid;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_2 <= __stream_conv2d_4_stream_ivalid_1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_3 <= __stream_conv2d_4_stream_ivalid_2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_4 <= __stream_conv2d_4_stream_ivalid_3;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_5 <= __stream_conv2d_4_stream_ivalid_4;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_6 <= __stream_conv2d_4_stream_ivalid_5;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_7 <= __stream_conv2d_4_stream_ivalid_6;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_8 <= __stream_conv2d_4_stream_ivalid_7;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_9 <= __stream_conv2d_4_stream_ivalid_8;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_10 <= __stream_conv2d_4_stream_ivalid_9;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_11 <= __stream_conv2d_4_stream_ivalid_10;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_12 <= __stream_conv2d_4_stream_ivalid_11;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_13 <= __stream_conv2d_4_stream_ivalid_12;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_14 <= __stream_conv2d_4_stream_ivalid_13;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_15 <= __stream_conv2d_4_stream_ivalid_14;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_16 <= __stream_conv2d_4_stream_ivalid_15;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_17 <= __stream_conv2d_4_stream_ivalid_16;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_18 <= __stream_conv2d_4_stream_ivalid_17;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_19 <= __stream_conv2d_4_stream_ivalid_18;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_20 <= __stream_conv2d_4_stream_ivalid_19;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_21 <= __stream_conv2d_4_stream_ivalid_20;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_22 <= __stream_conv2d_4_stream_ivalid_21;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_23 <= __stream_conv2d_4_stream_ivalid_22;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_24 <= __stream_conv2d_4_stream_ivalid_23;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_25 <= __stream_conv2d_4_stream_ivalid_24;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_26 <= __stream_conv2d_4_stream_ivalid_25;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_27 <= __stream_conv2d_4_stream_ivalid_26;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_28 <= __stream_conv2d_4_stream_ivalid_27;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_29 <= __stream_conv2d_4_stream_ivalid_28;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_30 <= __stream_conv2d_4_stream_ivalid_29;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_31 <= __stream_conv2d_4_stream_ivalid_30;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_402 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_406 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_409 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_412 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_416 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_419 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_422 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_426 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_429 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_432 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_436 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_439 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_442 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_446 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_449 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_452 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_456 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_459 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_462 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_466 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_469 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_472 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_476 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_479 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_482 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_486 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_489 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_492 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_496 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_499 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_502 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_506 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_509 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_512 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_516 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_519 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_522 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_526 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_529 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_532 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_536 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_539 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_542 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_546 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_549 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_552 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_556 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_559 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_562 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_566 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_569 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_572 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_576 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_579 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_734 <= _cond_data_374 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_753 <= _cond_data_374 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_772 <= _cond_data_374 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_791 <= _cond_data_374 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_810 <= _cond_data_374 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_829 <= _cond_data_374 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_848 <= _cond_data_374 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_867 <= _cond_data_374 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_886 <= _cond_data_374 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_902 <= _cond_data_381 + stream_conv2d_4_parameter_17_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_921 <= _cond_data_388 + stream_conv2d_4_parameter_18_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1254__variable_395 <= stream_conv2d_4_source_22_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1255__variable_394 <= stream_conv2d_4_source_21_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1256__variable_393 <= stream_conv2d_4_source_20_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1257__variable_398 <= stream_conv2d_4_source_25_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1258__variable_397 <= stream_conv2d_4_source_24_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1259__variable_396 <= stream_conv2d_4_source_23_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1260__variable_401 <= stream_conv2d_4_source_28_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1261__variable_400 <= stream_conv2d_4_source_27_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1262__variable_399 <= stream_conv2d_4_source_26_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1263_pointer_681 <= _pointer_data_681;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1264_reinterpretcast_672 <= _reinterpretcast_data_672;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1265_pointer_683 <= _pointer_data_683;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1266_reinterpretcast_673 <= _reinterpretcast_data_673;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1267_pointer_685 <= _pointer_data_685;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1268_reinterpretcast_674 <= _reinterpretcast_data_674;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1269_pointer_687 <= _pointer_data_687;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1270_reinterpretcast_675 <= _reinterpretcast_data_675;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1271_pointer_689 <= _pointer_data_689;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1272_reinterpretcast_676 <= _reinterpretcast_data_676;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1273_pointer_691 <= _pointer_data_691;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1274_reinterpretcast_677 <= _reinterpretcast_data_677;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1275_pointer_693 <= _pointer_data_693;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1276_reinterpretcast_678 <= _reinterpretcast_data_678;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1277_pointer_695 <= _pointer_data_695;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1278_reinterpretcast_679 <= _reinterpretcast_data_679;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1279_pointer_697 <= _pointer_data_697;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1280_reinterpretcast_680 <= _reinterpretcast_data_680;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1281__variable_344 <= stream_conv2d_4__reduce_reset_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1306__variable_339 <= stream_conv2d_4_parameter_0_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1319_cond_360 <= _cond_data_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1338_cond_367 <= _cond_data_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1282__delay_1281__variable_344 <= __delay_data_1281__variable_344;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1294_plus_902 <= _plus_data_902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1307__delay_1306__variable_339 <= __delay_data_1306__variable_339;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1320__delay_1319_cond_360 <= __delay_data_1319_cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1339__delay_1338_cond_367 <= __delay_data_1338_cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1358_plus_921 <= _plus_data_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1283__delay_1282__delay_1281__variable_344 <= __delay_data_1282__delay_1281__variable_344;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1295__delay_1294_plus_902 <= __delay_data_1294_plus_902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1308__delay_1307__delay_1306__variable_339 <= __delay_data_1307__delay_1306__variable_339;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1321__delay_1320__delay_1319_cond_360 <= __delay_data_1320__delay_1319_cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1340__delay_1339__delay_1338_cond_367 <= __delay_data_1339__delay_1338_cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1359__delay_1358_plus_921 <= __delay_data_1358_plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1284__delay_1283__delay_1282____variable_344 <= __delay_data_1283__delay_1282__delay_1281__variable_344;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1296__delay_1295__delay_1294_plus_902 <= __delay_data_1295__delay_1294_plus_902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1309__delay_1308__delay_1307____variable_339 <= __delay_data_1308__delay_1307__delay_1306__variable_339;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1322__delay_1321__delay_1320__delay_1319_cond_360 <= __delay_data_1321__delay_1320__delay_1319_cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1341__delay_1340__delay_1339__delay_1338_cond_367 <= __delay_data_1340__delay_1339__delay_1338_cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1360__delay_1359__delay_1358_plus_921 <= __delay_data_1359__delay_1358_plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1285__delay_1284__delay_1283____variable_344 <= __delay_data_1284__delay_1283__delay_1282____variable_344;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1297__delay_1296__delay_1295__delay_1294_plus_902 <= __delay_data_1296__delay_1295__delay_1294_plus_902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1310__delay_1309__delay_1308____variable_339 <= __delay_data_1309__delay_1308__delay_1307____variable_339;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1323__delay_1322__delay_1321__delay_1320___cond_360 <= __delay_data_1322__delay_1321__delay_1320__delay_1319_cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1342__delay_1341__delay_1340__delay_1339___cond_367 <= __delay_data_1341__delay_1340__delay_1339__delay_1338_cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1361__delay_1360__delay_1359__delay_1358_plus_921 <= __delay_data_1360__delay_1359__delay_1358_plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1286__delay_1285__delay_1284____variable_344 <= __delay_data_1285__delay_1284__delay_1283____variable_344;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1298__delay_1297__delay_1296__delay_1295___plus_902 <= __delay_data_1297__delay_1296__delay_1295__delay_1294_plus_902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1311__delay_1310__delay_1309____variable_339 <= __delay_data_1310__delay_1309__delay_1308____variable_339;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1324__delay_1323__delay_1322__delay_1321___cond_360 <= __delay_data_1323__delay_1322__delay_1321__delay_1320___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1343__delay_1342__delay_1341__delay_1340___cond_367 <= __delay_data_1342__delay_1341__delay_1340__delay_1339___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1362__delay_1361__delay_1360__delay_1359___plus_921 <= __delay_data_1361__delay_1360__delay_1359__delay_1358_plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1287__delay_1286__delay_1285____variable_344 <= __delay_data_1286__delay_1285__delay_1284____variable_344;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1299__delay_1298__delay_1297__delay_1296___plus_902 <= __delay_data_1298__delay_1297__delay_1296__delay_1295___plus_902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1312__delay_1311__delay_1310____variable_339 <= __delay_data_1311__delay_1310__delay_1309____variable_339;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1325__delay_1324__delay_1323__delay_1322___cond_360 <= __delay_data_1324__delay_1323__delay_1322__delay_1321___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1344__delay_1343__delay_1342__delay_1341___cond_367 <= __delay_data_1343__delay_1342__delay_1341__delay_1340___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1363__delay_1362__delay_1361__delay_1360___plus_921 <= __delay_data_1362__delay_1361__delay_1360__delay_1359___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1288__delay_1287__delay_1286____variable_344 <= __delay_data_1287__delay_1286__delay_1285____variable_344;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1300__delay_1299__delay_1298__delay_1297___plus_902 <= __delay_data_1299__delay_1298__delay_1297__delay_1296___plus_902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1313__delay_1312__delay_1311____variable_339 <= __delay_data_1312__delay_1311__delay_1310____variable_339;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1326__delay_1325__delay_1324__delay_1323___cond_360 <= __delay_data_1325__delay_1324__delay_1323__delay_1322___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1345__delay_1344__delay_1343__delay_1342___cond_367 <= __delay_data_1344__delay_1343__delay_1342__delay_1341___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1364__delay_1363__delay_1362__delay_1361___plus_921 <= __delay_data_1363__delay_1362__delay_1361__delay_1360___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1289__delay_1288__delay_1287____variable_344 <= __delay_data_1288__delay_1287__delay_1286____variable_344;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1301__delay_1300__delay_1299__delay_1298___plus_902 <= __delay_data_1300__delay_1299__delay_1298__delay_1297___plus_902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1314__delay_1313__delay_1312____variable_339 <= __delay_data_1313__delay_1312__delay_1311____variable_339;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1327__delay_1326__delay_1325__delay_1324___cond_360 <= __delay_data_1326__delay_1325__delay_1324__delay_1323___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1346__delay_1345__delay_1344__delay_1343___cond_367 <= __delay_data_1345__delay_1344__delay_1343__delay_1342___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1365__delay_1364__delay_1363__delay_1362___plus_921 <= __delay_data_1364__delay_1363__delay_1362__delay_1361___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1290__delay_1289__delay_1288____variable_344 <= __delay_data_1289__delay_1288__delay_1287____variable_344;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1302__delay_1301__delay_1300__delay_1299___plus_902 <= __delay_data_1301__delay_1300__delay_1299__delay_1298___plus_902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1315__delay_1314__delay_1313____variable_339 <= __delay_data_1314__delay_1313__delay_1312____variable_339;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1328__delay_1327__delay_1326__delay_1325___cond_360 <= __delay_data_1327__delay_1326__delay_1325__delay_1324___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1347__delay_1346__delay_1345__delay_1344___cond_367 <= __delay_data_1346__delay_1345__delay_1344__delay_1343___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1366__delay_1365__delay_1364__delay_1363___plus_921 <= __delay_data_1365__delay_1364__delay_1363__delay_1362___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1291__delay_1290__delay_1289____variable_344 <= __delay_data_1290__delay_1289__delay_1288____variable_344;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1303__delay_1302__delay_1301__delay_1300___plus_902 <= __delay_data_1302__delay_1301__delay_1300__delay_1299___plus_902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1316__delay_1315__delay_1314____variable_339 <= __delay_data_1315__delay_1314__delay_1313____variable_339;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1329__delay_1328__delay_1327__delay_1326___cond_360 <= __delay_data_1328__delay_1327__delay_1326__delay_1325___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1348__delay_1347__delay_1346__delay_1345___cond_367 <= __delay_data_1347__delay_1346__delay_1345__delay_1344___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1367__delay_1366__delay_1365__delay_1364___plus_921 <= __delay_data_1366__delay_1365__delay_1364__delay_1363___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1292__delay_1291__delay_1290____variable_344 <= __delay_data_1291__delay_1290__delay_1289____variable_344;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1304__delay_1303__delay_1302__delay_1301___plus_902 <= __delay_data_1303__delay_1302__delay_1301__delay_1300___plus_902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1317__delay_1316__delay_1315____variable_339 <= __delay_data_1316__delay_1315__delay_1314____variable_339;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1330__delay_1329__delay_1328__delay_1327___cond_360 <= __delay_data_1329__delay_1328__delay_1327__delay_1326___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1349__delay_1348__delay_1347__delay_1346___cond_367 <= __delay_data_1348__delay_1347__delay_1346__delay_1345___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1368__delay_1367__delay_1366__delay_1365___plus_921 <= __delay_data_1367__delay_1366__delay_1365__delay_1364___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1293__delay_1292__delay_1291____variable_344 <= __delay_data_1292__delay_1291__delay_1290____variable_344;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1305__delay_1304__delay_1303__delay_1302___plus_902 <= __delay_data_1304__delay_1303__delay_1302__delay_1301___plus_902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1318__delay_1317__delay_1316____variable_339 <= __delay_data_1317__delay_1316__delay_1315____variable_339;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1331__delay_1330__delay_1329__delay_1328___cond_360 <= __delay_data_1330__delay_1329__delay_1328__delay_1327___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1350__delay_1349__delay_1348__delay_1347___cond_367 <= __delay_data_1349__delay_1348__delay_1347__delay_1346___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1369__delay_1368__delay_1367__delay_1366___plus_921 <= __delay_data_1368__delay_1367__delay_1366__delay_1365___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1332__delay_1331__delay_1330__delay_1329___cond_360 <= __delay_data_1331__delay_1330__delay_1329__delay_1328___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1351__delay_1350__delay_1349__delay_1348___cond_367 <= __delay_data_1350__delay_1349__delay_1348__delay_1347___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1370__delay_1369__delay_1368__delay_1367___plus_921 <= __delay_data_1369__delay_1368__delay_1367__delay_1366___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1333__delay_1332__delay_1331__delay_1330___cond_360 <= __delay_data_1332__delay_1331__delay_1330__delay_1329___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1352__delay_1351__delay_1350__delay_1349___cond_367 <= __delay_data_1351__delay_1350__delay_1349__delay_1348___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1371__delay_1370__delay_1369__delay_1368___plus_921 <= __delay_data_1370__delay_1369__delay_1368__delay_1367___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1334__delay_1333__delay_1332__delay_1331___cond_360 <= __delay_data_1333__delay_1332__delay_1331__delay_1330___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1353__delay_1352__delay_1351__delay_1350___cond_367 <= __delay_data_1352__delay_1351__delay_1350__delay_1349___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1372__delay_1371__delay_1370__delay_1369___plus_921 <= __delay_data_1371__delay_1370__delay_1369__delay_1368___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1335__delay_1334__delay_1333__delay_1332___cond_360 <= __delay_data_1334__delay_1333__delay_1332__delay_1331___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1354__delay_1353__delay_1352__delay_1351___cond_367 <= __delay_data_1353__delay_1352__delay_1351__delay_1350___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1373__delay_1372__delay_1371__delay_1370___plus_921 <= __delay_data_1372__delay_1371__delay_1370__delay_1369___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1336__delay_1335__delay_1334__delay_1333___cond_360 <= __delay_data_1335__delay_1334__delay_1333__delay_1332___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1355__delay_1354__delay_1353__delay_1352___cond_367 <= __delay_data_1354__delay_1353__delay_1352__delay_1351___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1374__delay_1373__delay_1372__delay_1371___plus_921 <= __delay_data_1373__delay_1372__delay_1371__delay_1370___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1337__delay_1336__delay_1335__delay_1334___cond_360 <= __delay_data_1336__delay_1335__delay_1334__delay_1333___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1356__delay_1355__delay_1354__delay_1353___cond_367 <= __delay_data_1355__delay_1354__delay_1353__delay_1352___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1375__delay_1374__delay_1373__delay_1372___plus_921 <= __delay_data_1374__delay_1373__delay_1372__delay_1371___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_905 <= __substreamoutput_data_903 + __delay_data_1337__delay_1336__delay_1335__delay_1334___cond_360;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1357__delay_1356__delay_1355__delay_1354___cond_367 <= __delay_data_1356__delay_1355__delay_1354__delay_1353___cond_367;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1376__delay_1375__delay_1374__delay_1373___plus_921 <= __delay_data_1375__delay_1374__delay_1373__delay_1372___plus_921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1378__substreamoutput_904 <= __substreamoutput_data_904;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1379__delay_1378__substreamoutput_904 <= __delay_data_1378__substreamoutput_904;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1380__delay_1379__delay_1378__substreamoutput_904 <= __delay_data_1379__delay_1378__substreamoutput_904;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1381__delay_1380__delay_1379____substreamoutput_904 <= __delay_data_1380__delay_1379__delay_1378__substreamoutput_904;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1382__delay_1381__delay_1380____substreamoutput_904 <= __delay_data_1381__delay_1380__delay_1379____substreamoutput_904;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1383__delay_1382__delay_1381____substreamoutput_904 <= __delay_data_1382__delay_1381__delay_1380____substreamoutput_904;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1384__delay_1383__delay_1382____substreamoutput_904 <= __delay_data_1383__delay_1382__delay_1381____substreamoutput_904;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1385__delay_1384__delay_1383____substreamoutput_904 <= __delay_data_1384__delay_1383__delay_1382____substreamoutput_904;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1386__delay_1385__delay_1384____substreamoutput_904 <= __delay_data_1385__delay_1384__delay_1383____substreamoutput_904;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1387__delay_1386__delay_1385____substreamoutput_904 <= __delay_data_1386__delay_1385__delay_1384____substreamoutput_904;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _greaterthan_data_924 <= __substreamoutput_data_922 > 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1377__substreamoutput_922 <= __substreamoutput_data_922;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1388__delay_1387__delay_1386____substreamoutput_904 <= __delay_data_1387__delay_1386__delay_1385____substreamoutput_904;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _cond_data_926 <= (_greaterthan_data_924)? __delay_data_1377__substreamoutput_922 : 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_1389__delay_1388__delay_1387____substreamoutput_904 <= __delay_data_1388__delay_1387__delay_1386____substreamoutput_904;
      end 
      if(_set_flag_328) begin
        _stream_conv2d_4_parameter_0_next_parameter_data <= cparam_conv2d_4_stream_reduce_size;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_339 <= _stream_conv2d_4_parameter_0_next_parameter_data;
      end 
      if(_set_flag_329) begin
        _stream_conv2d_4_parameter_1_next_parameter_data <= conv2d_4_col_select;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_340 <= _stream_conv2d_4_parameter_1_next_parameter_data;
      end 
      if(_set_flag_330) begin
        _stream_conv2d_4_parameter_2_next_parameter_data <= conv2d_4_row_select_buf;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_341 <= _stream_conv2d_4_parameter_2_next_parameter_data;
      end 
      if(_set_flag_331) begin
        _stream_conv2d_4_parameter_3_next_parameter_data <= conv2d_4_stream_pad_masks;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_342 <= _stream_conv2d_4_parameter_3_next_parameter_data;
      end 
      if(_set_flag_332) begin
        _stream_conv2d_4_parameter_4_next_parameter_data <= cparam_conv2d_4_stream_omit_mask;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_343 <= _stream_conv2d_4_parameter_4_next_parameter_data;
      end 
      if(_set_flag_333) begin
        _stream_conv2d_4_parameter_6_next_parameter_data <= cparam_conv2d_4_bias_scala;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_354 <= _stream_conv2d_4_parameter_6_next_parameter_data;
      end 
      if(_set_flag_334) begin
        _stream_conv2d_4_source_7_source_mode <= 5'b10;
        _stream_conv2d_4_source_7_source_offset <= (cparam_conv2d_4_bias_num == 1)? 0 : conv2d_4_och_count_buf;
      end 
      if(_set_flag_334) begin
        _source_stream_conv2d_4_source_7_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_7_pat_stride_0 <= 0;
      end 
      if(_set_flag_334) begin
        _source_stream_conv2d_4_source_7_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_7_pat_stride_1 <= (cparam_conv2d_4_bias_num == 1)? 0 : 1;
      end 
      if(_set_flag_334) begin
        _source_stream_conv2d_4_source_7_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_7_pat_stride_2 <= 0;
      end 
      if(_set_flag_334) begin
        _source_stream_conv2d_4_source_7_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_7_pat_stride_3 <= 0;
      end 
      if(_set_flag_334) begin
        _stream_conv2d_4_source_7_source_sel <= 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_source_offset_buf <= _stream_conv2d_4_source_7_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_count_0 <= _source_stream_conv2d_4_source_7_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_count_1 <= _source_stream_conv2d_4_source_7_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_count_2 <= _source_stream_conv2d_4_source_7_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_count_3 <= _source_stream_conv2d_4_source_7_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_size_buf_0 <= _source_stream_conv2d_4_source_7_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_size_buf_1 <= _source_stream_conv2d_4_source_7_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_size_buf_2 <= _source_stream_conv2d_4_source_7_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_size_buf_3 <= _source_stream_conv2d_4_source_7_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_stride_buf_0 <= _source_stream_conv2d_4_source_7_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_stride_buf_1 <= _source_stream_conv2d_4_source_7_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_stride_buf_2 <= _source_stream_conv2d_4_source_7_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_stride_buf_3 <= _source_stream_conv2d_4_source_7_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_355 <= _stream_conv2d_4_source_7_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_idle <= 0;
        _stream_conv2d_4_source_7_source_ram_raddr <= _stream_conv2d_4_source_7_source_pat_all_offset;
        _stream_conv2d_4_source_7_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_0 <= _source_stream_conv2d_4_source_7_pat_cur_offset_0 + _source_stream_conv2d_4_source_7_pat_stride_buf_0;
        _source_stream_conv2d_4_source_7_pat_count_0 <= _source_stream_conv2d_4_source_7_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_4_source_7_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_7_pat_count_0 <= _source_stream_conv2d_4_source_7_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_4_source_7_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_1 <= _source_stream_conv2d_4_source_7_pat_cur_offset_1 + _source_stream_conv2d_4_source_7_pat_stride_buf_1;
        _source_stream_conv2d_4_source_7_pat_count_1 <= _source_stream_conv2d_4_source_7_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_7_pat_count_1 <= _source_stream_conv2d_4_source_7_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_2 <= _source_stream_conv2d_4_source_7_pat_cur_offset_2 + _source_stream_conv2d_4_source_7_pat_stride_buf_2;
        _source_stream_conv2d_4_source_7_pat_count_2 <= _source_stream_conv2d_4_source_7_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_7_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_7_pat_count_2 <= _source_stream_conv2d_4_source_7_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0) && (_source_stream_conv2d_4_source_7_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_3 <= _source_stream_conv2d_4_source_7_pat_cur_offset_3 + _source_stream_conv2d_4_source_7_pat_stride_buf_3;
        _source_stream_conv2d_4_source_7_pat_count_3 <= _source_stream_conv2d_4_source_7_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0) && (_source_stream_conv2d_4_source_7_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_7_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_7_pat_count_3 <= _source_stream_conv2d_4_source_7_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_source_ram_renable <= 0;
        _stream_conv2d_4_source_7_idle <= 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_source_ram_renable <= 0;
        _stream_conv2d_4_source_7_idle <= 1;
      end 
      if(_set_flag_343) begin
        _stream_conv2d_4_parameter_8_next_parameter_data <= cparam_conv2d_4_scale_scala;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_361 <= _stream_conv2d_4_parameter_8_next_parameter_data;
      end 
      if(_set_flag_344) begin
        _stream_conv2d_4_source_9_source_mode <= 5'b10;
        _stream_conv2d_4_source_9_source_offset <= (cparam_conv2d_4_scale_num == 1)? 0 : conv2d_4_och_count_buf;
      end 
      if(_set_flag_344) begin
        _source_stream_conv2d_4_source_9_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_9_pat_stride_0 <= 0;
      end 
      if(_set_flag_344) begin
        _source_stream_conv2d_4_source_9_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_9_pat_stride_1 <= (cparam_conv2d_4_scale_num == 1)? 0 : 1;
      end 
      if(_set_flag_344) begin
        _source_stream_conv2d_4_source_9_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_9_pat_stride_2 <= 0;
      end 
      if(_set_flag_344) begin
        _source_stream_conv2d_4_source_9_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_9_pat_stride_3 <= 0;
      end 
      if(_set_flag_344) begin
        _stream_conv2d_4_source_9_source_sel <= 2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_source_offset_buf <= _stream_conv2d_4_source_9_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_count_0 <= _source_stream_conv2d_4_source_9_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_count_1 <= _source_stream_conv2d_4_source_9_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_count_2 <= _source_stream_conv2d_4_source_9_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_count_3 <= _source_stream_conv2d_4_source_9_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_size_buf_0 <= _source_stream_conv2d_4_source_9_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_size_buf_1 <= _source_stream_conv2d_4_source_9_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_size_buf_2 <= _source_stream_conv2d_4_source_9_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_size_buf_3 <= _source_stream_conv2d_4_source_9_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_stride_buf_0 <= _source_stream_conv2d_4_source_9_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_stride_buf_1 <= _source_stream_conv2d_4_source_9_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_stride_buf_2 <= _source_stream_conv2d_4_source_9_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_stride_buf_3 <= _source_stream_conv2d_4_source_9_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_362 <= _stream_conv2d_4_source_9_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_idle <= 0;
        _stream_conv2d_4_source_9_source_ram_raddr <= _stream_conv2d_4_source_9_source_pat_all_offset;
        _stream_conv2d_4_source_9_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_0 <= _source_stream_conv2d_4_source_9_pat_cur_offset_0 + _source_stream_conv2d_4_source_9_pat_stride_buf_0;
        _source_stream_conv2d_4_source_9_pat_count_0 <= _source_stream_conv2d_4_source_9_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_4_source_9_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_9_pat_count_0 <= _source_stream_conv2d_4_source_9_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_4_source_9_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_1 <= _source_stream_conv2d_4_source_9_pat_cur_offset_1 + _source_stream_conv2d_4_source_9_pat_stride_buf_1;
        _source_stream_conv2d_4_source_9_pat_count_1 <= _source_stream_conv2d_4_source_9_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_9_pat_count_1 <= _source_stream_conv2d_4_source_9_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_2 <= _source_stream_conv2d_4_source_9_pat_cur_offset_2 + _source_stream_conv2d_4_source_9_pat_stride_buf_2;
        _source_stream_conv2d_4_source_9_pat_count_2 <= _source_stream_conv2d_4_source_9_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_9_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_9_pat_count_2 <= _source_stream_conv2d_4_source_9_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0) && (_source_stream_conv2d_4_source_9_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_3 <= _source_stream_conv2d_4_source_9_pat_cur_offset_3 + _source_stream_conv2d_4_source_9_pat_stride_buf_3;
        _source_stream_conv2d_4_source_9_pat_count_3 <= _source_stream_conv2d_4_source_9_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0) && (_source_stream_conv2d_4_source_9_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_9_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_9_pat_count_3 <= _source_stream_conv2d_4_source_9_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_source_ram_renable <= 0;
        _stream_conv2d_4_source_9_idle <= 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_source_ram_renable <= 0;
        _stream_conv2d_4_source_9_idle <= 1;
      end 
      if(_set_flag_353) begin
        _stream_conv2d_4_parameter_10_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_368 <= _stream_conv2d_4_parameter_10_next_parameter_data;
      end 
      if(_set_flag_354) begin
        _stream_conv2d_4_source_11_source_mode <= 5'b0;
        _stream_conv2d_4_source_11_source_empty_data <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_11_source_mode & 5'b0))) begin
        _stream_conv2d_4_source_11_idle <= 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_11_source_mode & 5'b0)) && _stream_conv2d_4_is_root) begin
        __variable_wdata_369 <= _stream_conv2d_4_source_11_source_empty_data;
      end 
      if(_set_flag_355) begin
        _stream_conv2d_4_parameter_12_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_375 <= _stream_conv2d_4_parameter_12_next_parameter_data;
      end 
      if(_set_flag_356) begin
        _stream_conv2d_4_source_13_source_mode <= 5'b0;
        _stream_conv2d_4_source_13_source_empty_data <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_13_source_mode & 5'b0))) begin
        _stream_conv2d_4_source_13_idle <= 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_13_source_mode & 5'b0)) && _stream_conv2d_4_is_root) begin
        __variable_wdata_376 <= _stream_conv2d_4_source_13_source_empty_data;
      end 
      if(_set_flag_357) begin
        _stream_conv2d_4_parameter_14_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_382 <= _stream_conv2d_4_parameter_14_next_parameter_data;
      end 
      if(_set_flag_358) begin
        _stream_conv2d_4_source_15_source_mode <= 5'b0;
        _stream_conv2d_4_source_15_source_empty_data <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_15_source_mode & 5'b0))) begin
        _stream_conv2d_4_source_15_idle <= 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_15_source_mode & 5'b0)) && _stream_conv2d_4_is_root) begin
        __variable_wdata_383 <= _stream_conv2d_4_source_15_source_empty_data;
      end 
      if(_set_flag_359) begin
        _stream_conv2d_4_parameter_16_next_parameter_data <= cparam_conv2d_4_cshamt_mul_value;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_389 <= _stream_conv2d_4_parameter_16_next_parameter_data;
      end 
      if(_set_flag_360) begin
        _stream_conv2d_4_parameter_17_next_parameter_data <= cparam_conv2d_4_cshamt_sum_value;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_390 <= _stream_conv2d_4_parameter_17_next_parameter_data;
      end 
      if(_set_flag_361) begin
        _stream_conv2d_4_parameter_18_next_parameter_data <= cparam_conv2d_4_cshamt_out_value;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_391 <= _stream_conv2d_4_parameter_18_next_parameter_data;
      end 
      if(_set_flag_362) begin
        _stream_conv2d_4_parameter_19_next_parameter_data <= cparam_conv2d_4_act_func_index;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_392 <= _stream_conv2d_4_parameter_19_next_parameter_data;
      end 
      if(_set_flag_363) begin
        _stream_conv2d_4_source_20_source_mode <= 5'b10;
        _stream_conv2d_4_source_20_source_offset <= conv2d_4_stream_act_local_0 + conv2d_4_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_363) begin
        _source_stream_conv2d_4_source_20_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_20_pat_stride_0 <= 1;
      end 
      if(_set_flag_363) begin
        _source_stream_conv2d_4_source_20_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_20_pat_stride_1 <= 0;
      end 
      if(_set_flag_363) begin
        _source_stream_conv2d_4_source_20_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_20_pat_stride_2 <= 0;
      end 
      if(_set_flag_363) begin
        _source_stream_conv2d_4_source_20_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_20_pat_stride_3 <= 0;
      end 
      if(_set_flag_363) begin
        _stream_conv2d_4_source_20_source_sel <= 3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_source_offset_buf <= _stream_conv2d_4_source_20_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_count_0 <= _source_stream_conv2d_4_source_20_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_count_1 <= _source_stream_conv2d_4_source_20_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_count_2 <= _source_stream_conv2d_4_source_20_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_count_3 <= _source_stream_conv2d_4_source_20_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_size_buf_0 <= _source_stream_conv2d_4_source_20_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_size_buf_1 <= _source_stream_conv2d_4_source_20_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_size_buf_2 <= _source_stream_conv2d_4_source_20_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_size_buf_3 <= _source_stream_conv2d_4_source_20_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_stride_buf_0 <= _source_stream_conv2d_4_source_20_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_stride_buf_1 <= _source_stream_conv2d_4_source_20_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_stride_buf_2 <= _source_stream_conv2d_4_source_20_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_stride_buf_3 <= _source_stream_conv2d_4_source_20_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_393 <= _stream_conv2d_4_source_20_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_idle <= 0;
        _stream_conv2d_4_source_20_source_ram_raddr <= _stream_conv2d_4_source_20_source_pat_all_offset;
        _stream_conv2d_4_source_20_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_0 <= _source_stream_conv2d_4_source_20_pat_cur_offset_0 + _source_stream_conv2d_4_source_20_pat_stride_buf_0;
        _source_stream_conv2d_4_source_20_pat_count_0 <= _source_stream_conv2d_4_source_20_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_4_source_20_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_20_pat_count_0 <= _source_stream_conv2d_4_source_20_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_4_source_20_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_1 <= _source_stream_conv2d_4_source_20_pat_cur_offset_1 + _source_stream_conv2d_4_source_20_pat_stride_buf_1;
        _source_stream_conv2d_4_source_20_pat_count_1 <= _source_stream_conv2d_4_source_20_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_20_pat_count_1 <= _source_stream_conv2d_4_source_20_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_2 <= _source_stream_conv2d_4_source_20_pat_cur_offset_2 + _source_stream_conv2d_4_source_20_pat_stride_buf_2;
        _source_stream_conv2d_4_source_20_pat_count_2 <= _source_stream_conv2d_4_source_20_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_20_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_20_pat_count_2 <= _source_stream_conv2d_4_source_20_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0) && (_source_stream_conv2d_4_source_20_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_3 <= _source_stream_conv2d_4_source_20_pat_cur_offset_3 + _source_stream_conv2d_4_source_20_pat_stride_buf_3;
        _source_stream_conv2d_4_source_20_pat_count_3 <= _source_stream_conv2d_4_source_20_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0) && (_source_stream_conv2d_4_source_20_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_20_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_20_pat_count_3 <= _source_stream_conv2d_4_source_20_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_source_ram_renable <= 0;
        _stream_conv2d_4_source_20_idle <= 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_source_ram_renable <= 0;
        _stream_conv2d_4_source_20_idle <= 1;
      end 
      if(_set_flag_372) begin
        _stream_conv2d_4_source_21_source_mode <= 5'b10;
        _stream_conv2d_4_source_21_source_offset <= conv2d_4_stream_act_local_1 + conv2d_4_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_372) begin
        _source_stream_conv2d_4_source_21_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_21_pat_stride_0 <= 1;
      end 
      if(_set_flag_372) begin
        _source_stream_conv2d_4_source_21_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_21_pat_stride_1 <= 0;
      end 
      if(_set_flag_372) begin
        _source_stream_conv2d_4_source_21_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_21_pat_stride_2 <= 0;
      end 
      if(_set_flag_372) begin
        _source_stream_conv2d_4_source_21_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_21_pat_stride_3 <= 0;
      end 
      if(_set_flag_372) begin
        _stream_conv2d_4_source_21_source_sel <= 4;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_source_offset_buf <= _stream_conv2d_4_source_21_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_count_0 <= _source_stream_conv2d_4_source_21_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_count_1 <= _source_stream_conv2d_4_source_21_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_count_2 <= _source_stream_conv2d_4_source_21_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_count_3 <= _source_stream_conv2d_4_source_21_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_size_buf_0 <= _source_stream_conv2d_4_source_21_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_size_buf_1 <= _source_stream_conv2d_4_source_21_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_size_buf_2 <= _source_stream_conv2d_4_source_21_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_size_buf_3 <= _source_stream_conv2d_4_source_21_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_stride_buf_0 <= _source_stream_conv2d_4_source_21_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_stride_buf_1 <= _source_stream_conv2d_4_source_21_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_stride_buf_2 <= _source_stream_conv2d_4_source_21_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_stride_buf_3 <= _source_stream_conv2d_4_source_21_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_394 <= _stream_conv2d_4_source_21_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_idle <= 0;
        _stream_conv2d_4_source_21_source_ram_raddr <= _stream_conv2d_4_source_21_source_pat_all_offset;
        _stream_conv2d_4_source_21_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_0 <= _source_stream_conv2d_4_source_21_pat_cur_offset_0 + _source_stream_conv2d_4_source_21_pat_stride_buf_0;
        _source_stream_conv2d_4_source_21_pat_count_0 <= _source_stream_conv2d_4_source_21_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_4_source_21_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_21_pat_count_0 <= _source_stream_conv2d_4_source_21_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_4_source_21_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_1 <= _source_stream_conv2d_4_source_21_pat_cur_offset_1 + _source_stream_conv2d_4_source_21_pat_stride_buf_1;
        _source_stream_conv2d_4_source_21_pat_count_1 <= _source_stream_conv2d_4_source_21_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_21_pat_count_1 <= _source_stream_conv2d_4_source_21_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_2 <= _source_stream_conv2d_4_source_21_pat_cur_offset_2 + _source_stream_conv2d_4_source_21_pat_stride_buf_2;
        _source_stream_conv2d_4_source_21_pat_count_2 <= _source_stream_conv2d_4_source_21_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_21_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_21_pat_count_2 <= _source_stream_conv2d_4_source_21_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0) && (_source_stream_conv2d_4_source_21_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_3 <= _source_stream_conv2d_4_source_21_pat_cur_offset_3 + _source_stream_conv2d_4_source_21_pat_stride_buf_3;
        _source_stream_conv2d_4_source_21_pat_count_3 <= _source_stream_conv2d_4_source_21_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0) && (_source_stream_conv2d_4_source_21_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_21_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_21_pat_count_3 <= _source_stream_conv2d_4_source_21_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_source_ram_renable <= 0;
        _stream_conv2d_4_source_21_idle <= 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_source_ram_renable <= 0;
        _stream_conv2d_4_source_21_idle <= 1;
      end 
      if(_set_flag_381) begin
        _stream_conv2d_4_source_22_source_mode <= 5'b10;
        _stream_conv2d_4_source_22_source_offset <= conv2d_4_stream_act_local_2 + conv2d_4_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_381) begin
        _source_stream_conv2d_4_source_22_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_22_pat_stride_0 <= 1;
      end 
      if(_set_flag_381) begin
        _source_stream_conv2d_4_source_22_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_22_pat_stride_1 <= 0;
      end 
      if(_set_flag_381) begin
        _source_stream_conv2d_4_source_22_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_22_pat_stride_2 <= 0;
      end 
      if(_set_flag_381) begin
        _source_stream_conv2d_4_source_22_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_22_pat_stride_3 <= 0;
      end 
      if(_set_flag_381) begin
        _stream_conv2d_4_source_22_source_sel <= 5;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_source_offset_buf <= _stream_conv2d_4_source_22_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_count_0 <= _source_stream_conv2d_4_source_22_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_count_1 <= _source_stream_conv2d_4_source_22_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_count_2 <= _source_stream_conv2d_4_source_22_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_count_3 <= _source_stream_conv2d_4_source_22_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_size_buf_0 <= _source_stream_conv2d_4_source_22_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_size_buf_1 <= _source_stream_conv2d_4_source_22_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_size_buf_2 <= _source_stream_conv2d_4_source_22_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_size_buf_3 <= _source_stream_conv2d_4_source_22_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_stride_buf_0 <= _source_stream_conv2d_4_source_22_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_stride_buf_1 <= _source_stream_conv2d_4_source_22_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_stride_buf_2 <= _source_stream_conv2d_4_source_22_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_stride_buf_3 <= _source_stream_conv2d_4_source_22_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_395 <= _stream_conv2d_4_source_22_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_idle <= 0;
        _stream_conv2d_4_source_22_source_ram_raddr <= _stream_conv2d_4_source_22_source_pat_all_offset;
        _stream_conv2d_4_source_22_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_0 <= _source_stream_conv2d_4_source_22_pat_cur_offset_0 + _source_stream_conv2d_4_source_22_pat_stride_buf_0;
        _source_stream_conv2d_4_source_22_pat_count_0 <= _source_stream_conv2d_4_source_22_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_4_source_22_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_22_pat_count_0 <= _source_stream_conv2d_4_source_22_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_4_source_22_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_1 <= _source_stream_conv2d_4_source_22_pat_cur_offset_1 + _source_stream_conv2d_4_source_22_pat_stride_buf_1;
        _source_stream_conv2d_4_source_22_pat_count_1 <= _source_stream_conv2d_4_source_22_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_22_pat_count_1 <= _source_stream_conv2d_4_source_22_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_2 <= _source_stream_conv2d_4_source_22_pat_cur_offset_2 + _source_stream_conv2d_4_source_22_pat_stride_buf_2;
        _source_stream_conv2d_4_source_22_pat_count_2 <= _source_stream_conv2d_4_source_22_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_22_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_22_pat_count_2 <= _source_stream_conv2d_4_source_22_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0) && (_source_stream_conv2d_4_source_22_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_3 <= _source_stream_conv2d_4_source_22_pat_cur_offset_3 + _source_stream_conv2d_4_source_22_pat_stride_buf_3;
        _source_stream_conv2d_4_source_22_pat_count_3 <= _source_stream_conv2d_4_source_22_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0) && (_source_stream_conv2d_4_source_22_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_22_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_22_pat_count_3 <= _source_stream_conv2d_4_source_22_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_source_ram_renable <= 0;
        _stream_conv2d_4_source_22_idle <= 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_source_ram_renable <= 0;
        _stream_conv2d_4_source_22_idle <= 1;
      end 
      if(_set_flag_390) begin
        _stream_conv2d_4_source_23_source_mode <= 5'b10;
        _stream_conv2d_4_source_23_source_offset <= conv2d_4_stream_act_local_3 + conv2d_4_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_390) begin
        _source_stream_conv2d_4_source_23_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_23_pat_stride_0 <= 1;
      end 
      if(_set_flag_390) begin
        _source_stream_conv2d_4_source_23_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_23_pat_stride_1 <= 0;
      end 
      if(_set_flag_390) begin
        _source_stream_conv2d_4_source_23_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_23_pat_stride_2 <= 0;
      end 
      if(_set_flag_390) begin
        _source_stream_conv2d_4_source_23_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_23_pat_stride_3 <= 0;
      end 
      if(_set_flag_390) begin
        _stream_conv2d_4_source_23_source_sel <= 6;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_source_offset_buf <= _stream_conv2d_4_source_23_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_count_0 <= _source_stream_conv2d_4_source_23_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_count_1 <= _source_stream_conv2d_4_source_23_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_count_2 <= _source_stream_conv2d_4_source_23_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_count_3 <= _source_stream_conv2d_4_source_23_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_size_buf_0 <= _source_stream_conv2d_4_source_23_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_size_buf_1 <= _source_stream_conv2d_4_source_23_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_size_buf_2 <= _source_stream_conv2d_4_source_23_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_size_buf_3 <= _source_stream_conv2d_4_source_23_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_stride_buf_0 <= _source_stream_conv2d_4_source_23_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_stride_buf_1 <= _source_stream_conv2d_4_source_23_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_stride_buf_2 <= _source_stream_conv2d_4_source_23_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_stride_buf_3 <= _source_stream_conv2d_4_source_23_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_396 <= _stream_conv2d_4_source_23_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_idle <= 0;
        _stream_conv2d_4_source_23_source_ram_raddr <= _stream_conv2d_4_source_23_source_pat_all_offset;
        _stream_conv2d_4_source_23_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_0 <= _source_stream_conv2d_4_source_23_pat_cur_offset_0 + _source_stream_conv2d_4_source_23_pat_stride_buf_0;
        _source_stream_conv2d_4_source_23_pat_count_0 <= _source_stream_conv2d_4_source_23_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_4_source_23_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_23_pat_count_0 <= _source_stream_conv2d_4_source_23_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_4_source_23_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_1 <= _source_stream_conv2d_4_source_23_pat_cur_offset_1 + _source_stream_conv2d_4_source_23_pat_stride_buf_1;
        _source_stream_conv2d_4_source_23_pat_count_1 <= _source_stream_conv2d_4_source_23_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_23_pat_count_1 <= _source_stream_conv2d_4_source_23_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_2 <= _source_stream_conv2d_4_source_23_pat_cur_offset_2 + _source_stream_conv2d_4_source_23_pat_stride_buf_2;
        _source_stream_conv2d_4_source_23_pat_count_2 <= _source_stream_conv2d_4_source_23_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_23_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_23_pat_count_2 <= _source_stream_conv2d_4_source_23_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0) && (_source_stream_conv2d_4_source_23_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_3 <= _source_stream_conv2d_4_source_23_pat_cur_offset_3 + _source_stream_conv2d_4_source_23_pat_stride_buf_3;
        _source_stream_conv2d_4_source_23_pat_count_3 <= _source_stream_conv2d_4_source_23_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0) && (_source_stream_conv2d_4_source_23_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_23_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_23_pat_count_3 <= _source_stream_conv2d_4_source_23_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_source_ram_renable <= 0;
        _stream_conv2d_4_source_23_idle <= 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_source_ram_renable <= 0;
        _stream_conv2d_4_source_23_idle <= 1;
      end 
      if(_set_flag_399) begin
        _stream_conv2d_4_source_24_source_mode <= 5'b10;
        _stream_conv2d_4_source_24_source_offset <= conv2d_4_stream_act_local_4 + conv2d_4_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_399) begin
        _source_stream_conv2d_4_source_24_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_24_pat_stride_0 <= 1;
      end 
      if(_set_flag_399) begin
        _source_stream_conv2d_4_source_24_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_24_pat_stride_1 <= 0;
      end 
      if(_set_flag_399) begin
        _source_stream_conv2d_4_source_24_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_24_pat_stride_2 <= 0;
      end 
      if(_set_flag_399) begin
        _source_stream_conv2d_4_source_24_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_24_pat_stride_3 <= 0;
      end 
      if(_set_flag_399) begin
        _stream_conv2d_4_source_24_source_sel <= 7;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_source_offset_buf <= _stream_conv2d_4_source_24_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_count_0 <= _source_stream_conv2d_4_source_24_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_count_1 <= _source_stream_conv2d_4_source_24_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_count_2 <= _source_stream_conv2d_4_source_24_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_count_3 <= _source_stream_conv2d_4_source_24_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_size_buf_0 <= _source_stream_conv2d_4_source_24_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_size_buf_1 <= _source_stream_conv2d_4_source_24_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_size_buf_2 <= _source_stream_conv2d_4_source_24_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_size_buf_3 <= _source_stream_conv2d_4_source_24_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_stride_buf_0 <= _source_stream_conv2d_4_source_24_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_stride_buf_1 <= _source_stream_conv2d_4_source_24_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_stride_buf_2 <= _source_stream_conv2d_4_source_24_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_stride_buf_3 <= _source_stream_conv2d_4_source_24_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_397 <= _stream_conv2d_4_source_24_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_idle <= 0;
        _stream_conv2d_4_source_24_source_ram_raddr <= _stream_conv2d_4_source_24_source_pat_all_offset;
        _stream_conv2d_4_source_24_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_0 <= _source_stream_conv2d_4_source_24_pat_cur_offset_0 + _source_stream_conv2d_4_source_24_pat_stride_buf_0;
        _source_stream_conv2d_4_source_24_pat_count_0 <= _source_stream_conv2d_4_source_24_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_4_source_24_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_24_pat_count_0 <= _source_stream_conv2d_4_source_24_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_4_source_24_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_1 <= _source_stream_conv2d_4_source_24_pat_cur_offset_1 + _source_stream_conv2d_4_source_24_pat_stride_buf_1;
        _source_stream_conv2d_4_source_24_pat_count_1 <= _source_stream_conv2d_4_source_24_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_24_pat_count_1 <= _source_stream_conv2d_4_source_24_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_2 <= _source_stream_conv2d_4_source_24_pat_cur_offset_2 + _source_stream_conv2d_4_source_24_pat_stride_buf_2;
        _source_stream_conv2d_4_source_24_pat_count_2 <= _source_stream_conv2d_4_source_24_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_24_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_24_pat_count_2 <= _source_stream_conv2d_4_source_24_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0) && (_source_stream_conv2d_4_source_24_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_3 <= _source_stream_conv2d_4_source_24_pat_cur_offset_3 + _source_stream_conv2d_4_source_24_pat_stride_buf_3;
        _source_stream_conv2d_4_source_24_pat_count_3 <= _source_stream_conv2d_4_source_24_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0) && (_source_stream_conv2d_4_source_24_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_24_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_24_pat_count_3 <= _source_stream_conv2d_4_source_24_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_source_ram_renable <= 0;
        _stream_conv2d_4_source_24_idle <= 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_source_ram_renable <= 0;
        _stream_conv2d_4_source_24_idle <= 1;
      end 
      if(_set_flag_408) begin
        _stream_conv2d_4_source_25_source_mode <= 5'b10;
        _stream_conv2d_4_source_25_source_offset <= conv2d_4_stream_act_local_5 + conv2d_4_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_408) begin
        _source_stream_conv2d_4_source_25_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_25_pat_stride_0 <= 1;
      end 
      if(_set_flag_408) begin
        _source_stream_conv2d_4_source_25_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_25_pat_stride_1 <= 0;
      end 
      if(_set_flag_408) begin
        _source_stream_conv2d_4_source_25_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_25_pat_stride_2 <= 0;
      end 
      if(_set_flag_408) begin
        _source_stream_conv2d_4_source_25_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_25_pat_stride_3 <= 0;
      end 
      if(_set_flag_408) begin
        _stream_conv2d_4_source_25_source_sel <= 8;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_source_offset_buf <= _stream_conv2d_4_source_25_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_count_0 <= _source_stream_conv2d_4_source_25_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_count_1 <= _source_stream_conv2d_4_source_25_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_count_2 <= _source_stream_conv2d_4_source_25_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_count_3 <= _source_stream_conv2d_4_source_25_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_size_buf_0 <= _source_stream_conv2d_4_source_25_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_size_buf_1 <= _source_stream_conv2d_4_source_25_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_size_buf_2 <= _source_stream_conv2d_4_source_25_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_size_buf_3 <= _source_stream_conv2d_4_source_25_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_stride_buf_0 <= _source_stream_conv2d_4_source_25_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_stride_buf_1 <= _source_stream_conv2d_4_source_25_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_stride_buf_2 <= _source_stream_conv2d_4_source_25_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_stride_buf_3 <= _source_stream_conv2d_4_source_25_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_398 <= _stream_conv2d_4_source_25_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_idle <= 0;
        _stream_conv2d_4_source_25_source_ram_raddr <= _stream_conv2d_4_source_25_source_pat_all_offset;
        _stream_conv2d_4_source_25_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_0 <= _source_stream_conv2d_4_source_25_pat_cur_offset_0 + _source_stream_conv2d_4_source_25_pat_stride_buf_0;
        _source_stream_conv2d_4_source_25_pat_count_0 <= _source_stream_conv2d_4_source_25_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_4_source_25_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_25_pat_count_0 <= _source_stream_conv2d_4_source_25_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_4_source_25_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_1 <= _source_stream_conv2d_4_source_25_pat_cur_offset_1 + _source_stream_conv2d_4_source_25_pat_stride_buf_1;
        _source_stream_conv2d_4_source_25_pat_count_1 <= _source_stream_conv2d_4_source_25_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_25_pat_count_1 <= _source_stream_conv2d_4_source_25_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_2 <= _source_stream_conv2d_4_source_25_pat_cur_offset_2 + _source_stream_conv2d_4_source_25_pat_stride_buf_2;
        _source_stream_conv2d_4_source_25_pat_count_2 <= _source_stream_conv2d_4_source_25_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_25_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_25_pat_count_2 <= _source_stream_conv2d_4_source_25_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0) && (_source_stream_conv2d_4_source_25_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_3 <= _source_stream_conv2d_4_source_25_pat_cur_offset_3 + _source_stream_conv2d_4_source_25_pat_stride_buf_3;
        _source_stream_conv2d_4_source_25_pat_count_3 <= _source_stream_conv2d_4_source_25_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0) && (_source_stream_conv2d_4_source_25_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_25_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_25_pat_count_3 <= _source_stream_conv2d_4_source_25_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_source_ram_renable <= 0;
        _stream_conv2d_4_source_25_idle <= 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_source_ram_renable <= 0;
        _stream_conv2d_4_source_25_idle <= 1;
      end 
      if(_set_flag_417) begin
        _stream_conv2d_4_source_26_source_mode <= 5'b10;
        _stream_conv2d_4_source_26_source_offset <= conv2d_4_stream_act_local_6 + conv2d_4_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_417) begin
        _source_stream_conv2d_4_source_26_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_26_pat_stride_0 <= 1;
      end 
      if(_set_flag_417) begin
        _source_stream_conv2d_4_source_26_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_26_pat_stride_1 <= 0;
      end 
      if(_set_flag_417) begin
        _source_stream_conv2d_4_source_26_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_26_pat_stride_2 <= 0;
      end 
      if(_set_flag_417) begin
        _source_stream_conv2d_4_source_26_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_26_pat_stride_3 <= 0;
      end 
      if(_set_flag_417) begin
        _stream_conv2d_4_source_26_source_sel <= 9;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_source_offset_buf <= _stream_conv2d_4_source_26_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_count_0 <= _source_stream_conv2d_4_source_26_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_count_1 <= _source_stream_conv2d_4_source_26_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_count_2 <= _source_stream_conv2d_4_source_26_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_count_3 <= _source_stream_conv2d_4_source_26_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_size_buf_0 <= _source_stream_conv2d_4_source_26_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_size_buf_1 <= _source_stream_conv2d_4_source_26_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_size_buf_2 <= _source_stream_conv2d_4_source_26_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_size_buf_3 <= _source_stream_conv2d_4_source_26_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_stride_buf_0 <= _source_stream_conv2d_4_source_26_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_stride_buf_1 <= _source_stream_conv2d_4_source_26_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_stride_buf_2 <= _source_stream_conv2d_4_source_26_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_stride_buf_3 <= _source_stream_conv2d_4_source_26_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_399 <= _stream_conv2d_4_source_26_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_idle <= 0;
        _stream_conv2d_4_source_26_source_ram_raddr <= _stream_conv2d_4_source_26_source_pat_all_offset;
        _stream_conv2d_4_source_26_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_0 <= _source_stream_conv2d_4_source_26_pat_cur_offset_0 + _source_stream_conv2d_4_source_26_pat_stride_buf_0;
        _source_stream_conv2d_4_source_26_pat_count_0 <= _source_stream_conv2d_4_source_26_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_4_source_26_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_26_pat_count_0 <= _source_stream_conv2d_4_source_26_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_4_source_26_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_1 <= _source_stream_conv2d_4_source_26_pat_cur_offset_1 + _source_stream_conv2d_4_source_26_pat_stride_buf_1;
        _source_stream_conv2d_4_source_26_pat_count_1 <= _source_stream_conv2d_4_source_26_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_26_pat_count_1 <= _source_stream_conv2d_4_source_26_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_2 <= _source_stream_conv2d_4_source_26_pat_cur_offset_2 + _source_stream_conv2d_4_source_26_pat_stride_buf_2;
        _source_stream_conv2d_4_source_26_pat_count_2 <= _source_stream_conv2d_4_source_26_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_26_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_26_pat_count_2 <= _source_stream_conv2d_4_source_26_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0) && (_source_stream_conv2d_4_source_26_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_3 <= _source_stream_conv2d_4_source_26_pat_cur_offset_3 + _source_stream_conv2d_4_source_26_pat_stride_buf_3;
        _source_stream_conv2d_4_source_26_pat_count_3 <= _source_stream_conv2d_4_source_26_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0) && (_source_stream_conv2d_4_source_26_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_26_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_26_pat_count_3 <= _source_stream_conv2d_4_source_26_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_source_ram_renable <= 0;
        _stream_conv2d_4_source_26_idle <= 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_source_ram_renable <= 0;
        _stream_conv2d_4_source_26_idle <= 1;
      end 
      if(_set_flag_426) begin
        _stream_conv2d_4_source_27_source_mode <= 5'b10;
        _stream_conv2d_4_source_27_source_offset <= conv2d_4_stream_act_local_7 + conv2d_4_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_426) begin
        _source_stream_conv2d_4_source_27_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_27_pat_stride_0 <= 1;
      end 
      if(_set_flag_426) begin
        _source_stream_conv2d_4_source_27_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_27_pat_stride_1 <= 0;
      end 
      if(_set_flag_426) begin
        _source_stream_conv2d_4_source_27_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_27_pat_stride_2 <= 0;
      end 
      if(_set_flag_426) begin
        _source_stream_conv2d_4_source_27_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_27_pat_stride_3 <= 0;
      end 
      if(_set_flag_426) begin
        _stream_conv2d_4_source_27_source_sel <= 10;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_source_offset_buf <= _stream_conv2d_4_source_27_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_count_0 <= _source_stream_conv2d_4_source_27_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_count_1 <= _source_stream_conv2d_4_source_27_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_count_2 <= _source_stream_conv2d_4_source_27_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_count_3 <= _source_stream_conv2d_4_source_27_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_size_buf_0 <= _source_stream_conv2d_4_source_27_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_size_buf_1 <= _source_stream_conv2d_4_source_27_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_size_buf_2 <= _source_stream_conv2d_4_source_27_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_size_buf_3 <= _source_stream_conv2d_4_source_27_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_stride_buf_0 <= _source_stream_conv2d_4_source_27_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_stride_buf_1 <= _source_stream_conv2d_4_source_27_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_stride_buf_2 <= _source_stream_conv2d_4_source_27_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_stride_buf_3 <= _source_stream_conv2d_4_source_27_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_400 <= _stream_conv2d_4_source_27_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_idle <= 0;
        _stream_conv2d_4_source_27_source_ram_raddr <= _stream_conv2d_4_source_27_source_pat_all_offset;
        _stream_conv2d_4_source_27_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_0 <= _source_stream_conv2d_4_source_27_pat_cur_offset_0 + _source_stream_conv2d_4_source_27_pat_stride_buf_0;
        _source_stream_conv2d_4_source_27_pat_count_0 <= _source_stream_conv2d_4_source_27_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_4_source_27_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_27_pat_count_0 <= _source_stream_conv2d_4_source_27_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_4_source_27_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_1 <= _source_stream_conv2d_4_source_27_pat_cur_offset_1 + _source_stream_conv2d_4_source_27_pat_stride_buf_1;
        _source_stream_conv2d_4_source_27_pat_count_1 <= _source_stream_conv2d_4_source_27_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_27_pat_count_1 <= _source_stream_conv2d_4_source_27_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_2 <= _source_stream_conv2d_4_source_27_pat_cur_offset_2 + _source_stream_conv2d_4_source_27_pat_stride_buf_2;
        _source_stream_conv2d_4_source_27_pat_count_2 <= _source_stream_conv2d_4_source_27_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_27_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_27_pat_count_2 <= _source_stream_conv2d_4_source_27_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0) && (_source_stream_conv2d_4_source_27_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_3 <= _source_stream_conv2d_4_source_27_pat_cur_offset_3 + _source_stream_conv2d_4_source_27_pat_stride_buf_3;
        _source_stream_conv2d_4_source_27_pat_count_3 <= _source_stream_conv2d_4_source_27_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0) && (_source_stream_conv2d_4_source_27_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_27_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_27_pat_count_3 <= _source_stream_conv2d_4_source_27_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_source_ram_renable <= 0;
        _stream_conv2d_4_source_27_idle <= 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_source_ram_renable <= 0;
        _stream_conv2d_4_source_27_idle <= 1;
      end 
      if(_set_flag_435) begin
        _stream_conv2d_4_source_28_source_mode <= 5'b10;
        _stream_conv2d_4_source_28_source_offset <= conv2d_4_stream_act_local_8 + conv2d_4_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_435) begin
        _source_stream_conv2d_4_source_28_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_28_pat_stride_0 <= 1;
      end 
      if(_set_flag_435) begin
        _source_stream_conv2d_4_source_28_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_28_pat_stride_1 <= 0;
      end 
      if(_set_flag_435) begin
        _source_stream_conv2d_4_source_28_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_28_pat_stride_2 <= 0;
      end 
      if(_set_flag_435) begin
        _source_stream_conv2d_4_source_28_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_28_pat_stride_3 <= 0;
      end 
      if(_set_flag_435) begin
        _stream_conv2d_4_source_28_source_sel <= 11;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_source_offset_buf <= _stream_conv2d_4_source_28_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_count_0 <= _source_stream_conv2d_4_source_28_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_count_1 <= _source_stream_conv2d_4_source_28_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_count_2 <= _source_stream_conv2d_4_source_28_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_count_3 <= _source_stream_conv2d_4_source_28_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_size_buf_0 <= _source_stream_conv2d_4_source_28_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_size_buf_1 <= _source_stream_conv2d_4_source_28_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_size_buf_2 <= _source_stream_conv2d_4_source_28_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_size_buf_3 <= _source_stream_conv2d_4_source_28_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_stride_buf_0 <= _source_stream_conv2d_4_source_28_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_stride_buf_1 <= _source_stream_conv2d_4_source_28_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_stride_buf_2 <= _source_stream_conv2d_4_source_28_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_stride_buf_3 <= _source_stream_conv2d_4_source_28_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_401 <= _stream_conv2d_4_source_28_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_idle <= 0;
        _stream_conv2d_4_source_28_source_ram_raddr <= _stream_conv2d_4_source_28_source_pat_all_offset;
        _stream_conv2d_4_source_28_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_0 <= _source_stream_conv2d_4_source_28_pat_cur_offset_0 + _source_stream_conv2d_4_source_28_pat_stride_buf_0;
        _source_stream_conv2d_4_source_28_pat_count_0 <= _source_stream_conv2d_4_source_28_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_4_source_28_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_28_pat_count_0 <= _source_stream_conv2d_4_source_28_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_4_source_28_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_1 <= _source_stream_conv2d_4_source_28_pat_cur_offset_1 + _source_stream_conv2d_4_source_28_pat_stride_buf_1;
        _source_stream_conv2d_4_source_28_pat_count_1 <= _source_stream_conv2d_4_source_28_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_28_pat_count_1 <= _source_stream_conv2d_4_source_28_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_2 <= _source_stream_conv2d_4_source_28_pat_cur_offset_2 + _source_stream_conv2d_4_source_28_pat_stride_buf_2;
        _source_stream_conv2d_4_source_28_pat_count_2 <= _source_stream_conv2d_4_source_28_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_28_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_28_pat_count_2 <= _source_stream_conv2d_4_source_28_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0) && (_source_stream_conv2d_4_source_28_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_3 <= _source_stream_conv2d_4_source_28_pat_cur_offset_3 + _source_stream_conv2d_4_source_28_pat_stride_buf_3;
        _source_stream_conv2d_4_source_28_pat_count_3 <= _source_stream_conv2d_4_source_28_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0) && (_source_stream_conv2d_4_source_28_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_28_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_28_pat_count_3 <= _source_stream_conv2d_4_source_28_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_source_ram_renable <= 0;
        _stream_conv2d_4_source_28_idle <= 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_source_ram_renable <= 0;
        _stream_conv2d_4_source_28_idle <= 1;
      end 
      if(_set_flag_444) begin
        _stream_conv2d_4_source_29_source_mode <= 5'b10;
        _stream_conv2d_4_source_29_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_444) begin
        _source_stream_conv2d_4_source_29_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_29_pat_stride_0 <= 1;
      end 
      if(_set_flag_444) begin
        _source_stream_conv2d_4_source_29_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_29_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_444) begin
        _source_stream_conv2d_4_source_29_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_29_pat_stride_2 <= 0;
      end 
      if(_set_flag_444) begin
        _source_stream_conv2d_4_source_29_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_29_pat_stride_3 <= 0;
      end 
      if(_set_flag_444) begin
        _stream_conv2d_4_source_29_source_sel <= 12;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_source_offset_buf <= _stream_conv2d_4_source_29_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_count_0 <= _source_stream_conv2d_4_source_29_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_count_1 <= _source_stream_conv2d_4_source_29_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_count_2 <= _source_stream_conv2d_4_source_29_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_count_3 <= _source_stream_conv2d_4_source_29_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_size_buf_0 <= _source_stream_conv2d_4_source_29_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_size_buf_1 <= _source_stream_conv2d_4_source_29_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_size_buf_2 <= _source_stream_conv2d_4_source_29_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_size_buf_3 <= _source_stream_conv2d_4_source_29_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_stride_buf_0 <= _source_stream_conv2d_4_source_29_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_stride_buf_1 <= _source_stream_conv2d_4_source_29_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_stride_buf_2 <= _source_stream_conv2d_4_source_29_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_stride_buf_3 <= _source_stream_conv2d_4_source_29_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_627 <= _stream_conv2d_4_source_29_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_idle <= 0;
        _stream_conv2d_4_source_29_source_ram_raddr <= _stream_conv2d_4_source_29_source_pat_all_offset;
        _stream_conv2d_4_source_29_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_0 <= _source_stream_conv2d_4_source_29_pat_cur_offset_0 + _source_stream_conv2d_4_source_29_pat_stride_buf_0;
        _source_stream_conv2d_4_source_29_pat_count_0 <= _source_stream_conv2d_4_source_29_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_4_source_29_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_29_pat_count_0 <= _source_stream_conv2d_4_source_29_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_4_source_29_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_1 <= _source_stream_conv2d_4_source_29_pat_cur_offset_1 + _source_stream_conv2d_4_source_29_pat_stride_buf_1;
        _source_stream_conv2d_4_source_29_pat_count_1 <= _source_stream_conv2d_4_source_29_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_29_pat_count_1 <= _source_stream_conv2d_4_source_29_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_2 <= _source_stream_conv2d_4_source_29_pat_cur_offset_2 + _source_stream_conv2d_4_source_29_pat_stride_buf_2;
        _source_stream_conv2d_4_source_29_pat_count_2 <= _source_stream_conv2d_4_source_29_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_29_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_29_pat_count_2 <= _source_stream_conv2d_4_source_29_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0) && (_source_stream_conv2d_4_source_29_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_3 <= _source_stream_conv2d_4_source_29_pat_cur_offset_3 + _source_stream_conv2d_4_source_29_pat_stride_buf_3;
        _source_stream_conv2d_4_source_29_pat_count_3 <= _source_stream_conv2d_4_source_29_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0) && (_source_stream_conv2d_4_source_29_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_29_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_29_pat_count_3 <= _source_stream_conv2d_4_source_29_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_source_ram_renable <= 0;
        _stream_conv2d_4_source_29_idle <= 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_source_ram_renable <= 0;
        _stream_conv2d_4_source_29_idle <= 1;
      end 
      if(_set_flag_453) begin
        _stream_conv2d_4_source_30_source_mode <= 5'b10;
        _stream_conv2d_4_source_30_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_453) begin
        _source_stream_conv2d_4_source_30_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_30_pat_stride_0 <= 1;
      end 
      if(_set_flag_453) begin
        _source_stream_conv2d_4_source_30_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_30_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_453) begin
        _source_stream_conv2d_4_source_30_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_30_pat_stride_2 <= 0;
      end 
      if(_set_flag_453) begin
        _source_stream_conv2d_4_source_30_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_30_pat_stride_3 <= 0;
      end 
      if(_set_flag_453) begin
        _stream_conv2d_4_source_30_source_sel <= 13;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_source_offset_buf <= _stream_conv2d_4_source_30_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_count_0 <= _source_stream_conv2d_4_source_30_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_count_1 <= _source_stream_conv2d_4_source_30_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_count_2 <= _source_stream_conv2d_4_source_30_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_count_3 <= _source_stream_conv2d_4_source_30_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_size_buf_0 <= _source_stream_conv2d_4_source_30_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_size_buf_1 <= _source_stream_conv2d_4_source_30_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_size_buf_2 <= _source_stream_conv2d_4_source_30_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_size_buf_3 <= _source_stream_conv2d_4_source_30_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_stride_buf_0 <= _source_stream_conv2d_4_source_30_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_stride_buf_1 <= _source_stream_conv2d_4_source_30_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_stride_buf_2 <= _source_stream_conv2d_4_source_30_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_stride_buf_3 <= _source_stream_conv2d_4_source_30_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_628 <= _stream_conv2d_4_source_30_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_idle <= 0;
        _stream_conv2d_4_source_30_source_ram_raddr <= _stream_conv2d_4_source_30_source_pat_all_offset;
        _stream_conv2d_4_source_30_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_0 <= _source_stream_conv2d_4_source_30_pat_cur_offset_0 + _source_stream_conv2d_4_source_30_pat_stride_buf_0;
        _source_stream_conv2d_4_source_30_pat_count_0 <= _source_stream_conv2d_4_source_30_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_4_source_30_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_30_pat_count_0 <= _source_stream_conv2d_4_source_30_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_4_source_30_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_1 <= _source_stream_conv2d_4_source_30_pat_cur_offset_1 + _source_stream_conv2d_4_source_30_pat_stride_buf_1;
        _source_stream_conv2d_4_source_30_pat_count_1 <= _source_stream_conv2d_4_source_30_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_30_pat_count_1 <= _source_stream_conv2d_4_source_30_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_2 <= _source_stream_conv2d_4_source_30_pat_cur_offset_2 + _source_stream_conv2d_4_source_30_pat_stride_buf_2;
        _source_stream_conv2d_4_source_30_pat_count_2 <= _source_stream_conv2d_4_source_30_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_30_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_30_pat_count_2 <= _source_stream_conv2d_4_source_30_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0) && (_source_stream_conv2d_4_source_30_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_3 <= _source_stream_conv2d_4_source_30_pat_cur_offset_3 + _source_stream_conv2d_4_source_30_pat_stride_buf_3;
        _source_stream_conv2d_4_source_30_pat_count_3 <= _source_stream_conv2d_4_source_30_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0) && (_source_stream_conv2d_4_source_30_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_30_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_30_pat_count_3 <= _source_stream_conv2d_4_source_30_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_source_ram_renable <= 0;
        _stream_conv2d_4_source_30_idle <= 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_source_ram_renable <= 0;
        _stream_conv2d_4_source_30_idle <= 1;
      end 
      if(_set_flag_462) begin
        _stream_conv2d_4_source_31_source_mode <= 5'b10;
        _stream_conv2d_4_source_31_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_462) begin
        _source_stream_conv2d_4_source_31_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_31_pat_stride_0 <= 1;
      end 
      if(_set_flag_462) begin
        _source_stream_conv2d_4_source_31_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_31_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_462) begin
        _source_stream_conv2d_4_source_31_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_31_pat_stride_2 <= 0;
      end 
      if(_set_flag_462) begin
        _source_stream_conv2d_4_source_31_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_31_pat_stride_3 <= 0;
      end 
      if(_set_flag_462) begin
        _stream_conv2d_4_source_31_source_sel <= 14;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_source_offset_buf <= _stream_conv2d_4_source_31_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_count_0 <= _source_stream_conv2d_4_source_31_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_count_1 <= _source_stream_conv2d_4_source_31_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_count_2 <= _source_stream_conv2d_4_source_31_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_count_3 <= _source_stream_conv2d_4_source_31_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_size_buf_0 <= _source_stream_conv2d_4_source_31_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_size_buf_1 <= _source_stream_conv2d_4_source_31_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_size_buf_2 <= _source_stream_conv2d_4_source_31_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_size_buf_3 <= _source_stream_conv2d_4_source_31_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_stride_buf_0 <= _source_stream_conv2d_4_source_31_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_stride_buf_1 <= _source_stream_conv2d_4_source_31_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_stride_buf_2 <= _source_stream_conv2d_4_source_31_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_stride_buf_3 <= _source_stream_conv2d_4_source_31_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_629 <= _stream_conv2d_4_source_31_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_idle <= 0;
        _stream_conv2d_4_source_31_source_ram_raddr <= _stream_conv2d_4_source_31_source_pat_all_offset;
        _stream_conv2d_4_source_31_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_0 <= _source_stream_conv2d_4_source_31_pat_cur_offset_0 + _source_stream_conv2d_4_source_31_pat_stride_buf_0;
        _source_stream_conv2d_4_source_31_pat_count_0 <= _source_stream_conv2d_4_source_31_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_4_source_31_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_31_pat_count_0 <= _source_stream_conv2d_4_source_31_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_4_source_31_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_1 <= _source_stream_conv2d_4_source_31_pat_cur_offset_1 + _source_stream_conv2d_4_source_31_pat_stride_buf_1;
        _source_stream_conv2d_4_source_31_pat_count_1 <= _source_stream_conv2d_4_source_31_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_31_pat_count_1 <= _source_stream_conv2d_4_source_31_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_2 <= _source_stream_conv2d_4_source_31_pat_cur_offset_2 + _source_stream_conv2d_4_source_31_pat_stride_buf_2;
        _source_stream_conv2d_4_source_31_pat_count_2 <= _source_stream_conv2d_4_source_31_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_31_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_31_pat_count_2 <= _source_stream_conv2d_4_source_31_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0) && (_source_stream_conv2d_4_source_31_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_3 <= _source_stream_conv2d_4_source_31_pat_cur_offset_3 + _source_stream_conv2d_4_source_31_pat_stride_buf_3;
        _source_stream_conv2d_4_source_31_pat_count_3 <= _source_stream_conv2d_4_source_31_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0) && (_source_stream_conv2d_4_source_31_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_31_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_31_pat_count_3 <= _source_stream_conv2d_4_source_31_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_source_ram_renable <= 0;
        _stream_conv2d_4_source_31_idle <= 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_source_ram_renable <= 0;
        _stream_conv2d_4_source_31_idle <= 1;
      end 
      if(_set_flag_471) begin
        _stream_conv2d_4_source_32_source_mode <= 5'b10;
        _stream_conv2d_4_source_32_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_471) begin
        _source_stream_conv2d_4_source_32_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_32_pat_stride_0 <= 1;
      end 
      if(_set_flag_471) begin
        _source_stream_conv2d_4_source_32_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_32_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_471) begin
        _source_stream_conv2d_4_source_32_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_32_pat_stride_2 <= 0;
      end 
      if(_set_flag_471) begin
        _source_stream_conv2d_4_source_32_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_32_pat_stride_3 <= 0;
      end 
      if(_set_flag_471) begin
        _stream_conv2d_4_source_32_source_sel <= 15;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_source_offset_buf <= _stream_conv2d_4_source_32_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_count_0 <= _source_stream_conv2d_4_source_32_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_count_1 <= _source_stream_conv2d_4_source_32_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_count_2 <= _source_stream_conv2d_4_source_32_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_count_3 <= _source_stream_conv2d_4_source_32_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_size_buf_0 <= _source_stream_conv2d_4_source_32_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_size_buf_1 <= _source_stream_conv2d_4_source_32_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_size_buf_2 <= _source_stream_conv2d_4_source_32_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_size_buf_3 <= _source_stream_conv2d_4_source_32_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_stride_buf_0 <= _source_stream_conv2d_4_source_32_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_stride_buf_1 <= _source_stream_conv2d_4_source_32_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_stride_buf_2 <= _source_stream_conv2d_4_source_32_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_stride_buf_3 <= _source_stream_conv2d_4_source_32_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_630 <= _stream_conv2d_4_source_32_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_idle <= 0;
        _stream_conv2d_4_source_32_source_ram_raddr <= _stream_conv2d_4_source_32_source_pat_all_offset;
        _stream_conv2d_4_source_32_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_0 <= _source_stream_conv2d_4_source_32_pat_cur_offset_0 + _source_stream_conv2d_4_source_32_pat_stride_buf_0;
        _source_stream_conv2d_4_source_32_pat_count_0 <= _source_stream_conv2d_4_source_32_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_4_source_32_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_32_pat_count_0 <= _source_stream_conv2d_4_source_32_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_4_source_32_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_1 <= _source_stream_conv2d_4_source_32_pat_cur_offset_1 + _source_stream_conv2d_4_source_32_pat_stride_buf_1;
        _source_stream_conv2d_4_source_32_pat_count_1 <= _source_stream_conv2d_4_source_32_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_32_pat_count_1 <= _source_stream_conv2d_4_source_32_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_2 <= _source_stream_conv2d_4_source_32_pat_cur_offset_2 + _source_stream_conv2d_4_source_32_pat_stride_buf_2;
        _source_stream_conv2d_4_source_32_pat_count_2 <= _source_stream_conv2d_4_source_32_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_32_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_32_pat_count_2 <= _source_stream_conv2d_4_source_32_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0) && (_source_stream_conv2d_4_source_32_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_3 <= _source_stream_conv2d_4_source_32_pat_cur_offset_3 + _source_stream_conv2d_4_source_32_pat_stride_buf_3;
        _source_stream_conv2d_4_source_32_pat_count_3 <= _source_stream_conv2d_4_source_32_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0) && (_source_stream_conv2d_4_source_32_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_32_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_32_pat_count_3 <= _source_stream_conv2d_4_source_32_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_source_ram_renable <= 0;
        _stream_conv2d_4_source_32_idle <= 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_source_ram_renable <= 0;
        _stream_conv2d_4_source_32_idle <= 1;
      end 
      if(_set_flag_480) begin
        _stream_conv2d_4_source_33_source_mode <= 5'b10;
        _stream_conv2d_4_source_33_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_480) begin
        _source_stream_conv2d_4_source_33_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_33_pat_stride_0 <= 1;
      end 
      if(_set_flag_480) begin
        _source_stream_conv2d_4_source_33_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_33_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_480) begin
        _source_stream_conv2d_4_source_33_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_33_pat_stride_2 <= 0;
      end 
      if(_set_flag_480) begin
        _source_stream_conv2d_4_source_33_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_33_pat_stride_3 <= 0;
      end 
      if(_set_flag_480) begin
        _stream_conv2d_4_source_33_source_sel <= 16;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_source_offset_buf <= _stream_conv2d_4_source_33_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_count_0 <= _source_stream_conv2d_4_source_33_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_count_1 <= _source_stream_conv2d_4_source_33_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_count_2 <= _source_stream_conv2d_4_source_33_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_count_3 <= _source_stream_conv2d_4_source_33_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_size_buf_0 <= _source_stream_conv2d_4_source_33_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_size_buf_1 <= _source_stream_conv2d_4_source_33_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_size_buf_2 <= _source_stream_conv2d_4_source_33_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_size_buf_3 <= _source_stream_conv2d_4_source_33_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_stride_buf_0 <= _source_stream_conv2d_4_source_33_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_stride_buf_1 <= _source_stream_conv2d_4_source_33_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_stride_buf_2 <= _source_stream_conv2d_4_source_33_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_stride_buf_3 <= _source_stream_conv2d_4_source_33_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_631 <= _stream_conv2d_4_source_33_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_idle <= 0;
        _stream_conv2d_4_source_33_source_ram_raddr <= _stream_conv2d_4_source_33_source_pat_all_offset;
        _stream_conv2d_4_source_33_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_0 <= _source_stream_conv2d_4_source_33_pat_cur_offset_0 + _source_stream_conv2d_4_source_33_pat_stride_buf_0;
        _source_stream_conv2d_4_source_33_pat_count_0 <= _source_stream_conv2d_4_source_33_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_4_source_33_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_33_pat_count_0 <= _source_stream_conv2d_4_source_33_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_4_source_33_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_1 <= _source_stream_conv2d_4_source_33_pat_cur_offset_1 + _source_stream_conv2d_4_source_33_pat_stride_buf_1;
        _source_stream_conv2d_4_source_33_pat_count_1 <= _source_stream_conv2d_4_source_33_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_33_pat_count_1 <= _source_stream_conv2d_4_source_33_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_2 <= _source_stream_conv2d_4_source_33_pat_cur_offset_2 + _source_stream_conv2d_4_source_33_pat_stride_buf_2;
        _source_stream_conv2d_4_source_33_pat_count_2 <= _source_stream_conv2d_4_source_33_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_33_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_33_pat_count_2 <= _source_stream_conv2d_4_source_33_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0) && (_source_stream_conv2d_4_source_33_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_3 <= _source_stream_conv2d_4_source_33_pat_cur_offset_3 + _source_stream_conv2d_4_source_33_pat_stride_buf_3;
        _source_stream_conv2d_4_source_33_pat_count_3 <= _source_stream_conv2d_4_source_33_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0) && (_source_stream_conv2d_4_source_33_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_33_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_33_pat_count_3 <= _source_stream_conv2d_4_source_33_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_source_ram_renable <= 0;
        _stream_conv2d_4_source_33_idle <= 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_source_ram_renable <= 0;
        _stream_conv2d_4_source_33_idle <= 1;
      end 
      if(_set_flag_489) begin
        _stream_conv2d_4_source_34_source_mode <= 5'b10;
        _stream_conv2d_4_source_34_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_489) begin
        _source_stream_conv2d_4_source_34_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_34_pat_stride_0 <= 1;
      end 
      if(_set_flag_489) begin
        _source_stream_conv2d_4_source_34_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_34_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_489) begin
        _source_stream_conv2d_4_source_34_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_34_pat_stride_2 <= 0;
      end 
      if(_set_flag_489) begin
        _source_stream_conv2d_4_source_34_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_34_pat_stride_3 <= 0;
      end 
      if(_set_flag_489) begin
        _stream_conv2d_4_source_34_source_sel <= 17;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_source_offset_buf <= _stream_conv2d_4_source_34_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_count_0 <= _source_stream_conv2d_4_source_34_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_count_1 <= _source_stream_conv2d_4_source_34_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_count_2 <= _source_stream_conv2d_4_source_34_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_count_3 <= _source_stream_conv2d_4_source_34_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_size_buf_0 <= _source_stream_conv2d_4_source_34_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_size_buf_1 <= _source_stream_conv2d_4_source_34_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_size_buf_2 <= _source_stream_conv2d_4_source_34_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_size_buf_3 <= _source_stream_conv2d_4_source_34_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_stride_buf_0 <= _source_stream_conv2d_4_source_34_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_stride_buf_1 <= _source_stream_conv2d_4_source_34_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_stride_buf_2 <= _source_stream_conv2d_4_source_34_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_stride_buf_3 <= _source_stream_conv2d_4_source_34_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_632 <= _stream_conv2d_4_source_34_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_idle <= 0;
        _stream_conv2d_4_source_34_source_ram_raddr <= _stream_conv2d_4_source_34_source_pat_all_offset;
        _stream_conv2d_4_source_34_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_0 <= _source_stream_conv2d_4_source_34_pat_cur_offset_0 + _source_stream_conv2d_4_source_34_pat_stride_buf_0;
        _source_stream_conv2d_4_source_34_pat_count_0 <= _source_stream_conv2d_4_source_34_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_4_source_34_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_34_pat_count_0 <= _source_stream_conv2d_4_source_34_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_4_source_34_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_1 <= _source_stream_conv2d_4_source_34_pat_cur_offset_1 + _source_stream_conv2d_4_source_34_pat_stride_buf_1;
        _source_stream_conv2d_4_source_34_pat_count_1 <= _source_stream_conv2d_4_source_34_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_34_pat_count_1 <= _source_stream_conv2d_4_source_34_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_2 <= _source_stream_conv2d_4_source_34_pat_cur_offset_2 + _source_stream_conv2d_4_source_34_pat_stride_buf_2;
        _source_stream_conv2d_4_source_34_pat_count_2 <= _source_stream_conv2d_4_source_34_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_34_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_34_pat_count_2 <= _source_stream_conv2d_4_source_34_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0) && (_source_stream_conv2d_4_source_34_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_3 <= _source_stream_conv2d_4_source_34_pat_cur_offset_3 + _source_stream_conv2d_4_source_34_pat_stride_buf_3;
        _source_stream_conv2d_4_source_34_pat_count_3 <= _source_stream_conv2d_4_source_34_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0) && (_source_stream_conv2d_4_source_34_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_34_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_34_pat_count_3 <= _source_stream_conv2d_4_source_34_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_source_ram_renable <= 0;
        _stream_conv2d_4_source_34_idle <= 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_source_ram_renable <= 0;
        _stream_conv2d_4_source_34_idle <= 1;
      end 
      if(_set_flag_498) begin
        _stream_conv2d_4_source_35_source_mode <= 5'b10;
        _stream_conv2d_4_source_35_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_498) begin
        _source_stream_conv2d_4_source_35_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_35_pat_stride_0 <= 1;
      end 
      if(_set_flag_498) begin
        _source_stream_conv2d_4_source_35_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_35_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_498) begin
        _source_stream_conv2d_4_source_35_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_35_pat_stride_2 <= 0;
      end 
      if(_set_flag_498) begin
        _source_stream_conv2d_4_source_35_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_35_pat_stride_3 <= 0;
      end 
      if(_set_flag_498) begin
        _stream_conv2d_4_source_35_source_sel <= 18;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_source_offset_buf <= _stream_conv2d_4_source_35_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_count_0 <= _source_stream_conv2d_4_source_35_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_count_1 <= _source_stream_conv2d_4_source_35_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_count_2 <= _source_stream_conv2d_4_source_35_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_count_3 <= _source_stream_conv2d_4_source_35_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_size_buf_0 <= _source_stream_conv2d_4_source_35_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_size_buf_1 <= _source_stream_conv2d_4_source_35_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_size_buf_2 <= _source_stream_conv2d_4_source_35_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_size_buf_3 <= _source_stream_conv2d_4_source_35_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_stride_buf_0 <= _source_stream_conv2d_4_source_35_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_stride_buf_1 <= _source_stream_conv2d_4_source_35_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_stride_buf_2 <= _source_stream_conv2d_4_source_35_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_stride_buf_3 <= _source_stream_conv2d_4_source_35_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_633 <= _stream_conv2d_4_source_35_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_idle <= 0;
        _stream_conv2d_4_source_35_source_ram_raddr <= _stream_conv2d_4_source_35_source_pat_all_offset;
        _stream_conv2d_4_source_35_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_0 <= _source_stream_conv2d_4_source_35_pat_cur_offset_0 + _source_stream_conv2d_4_source_35_pat_stride_buf_0;
        _source_stream_conv2d_4_source_35_pat_count_0 <= _source_stream_conv2d_4_source_35_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_4_source_35_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_35_pat_count_0 <= _source_stream_conv2d_4_source_35_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_4_source_35_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_1 <= _source_stream_conv2d_4_source_35_pat_cur_offset_1 + _source_stream_conv2d_4_source_35_pat_stride_buf_1;
        _source_stream_conv2d_4_source_35_pat_count_1 <= _source_stream_conv2d_4_source_35_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_35_pat_count_1 <= _source_stream_conv2d_4_source_35_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_2 <= _source_stream_conv2d_4_source_35_pat_cur_offset_2 + _source_stream_conv2d_4_source_35_pat_stride_buf_2;
        _source_stream_conv2d_4_source_35_pat_count_2 <= _source_stream_conv2d_4_source_35_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_35_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_35_pat_count_2 <= _source_stream_conv2d_4_source_35_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0) && (_source_stream_conv2d_4_source_35_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_3 <= _source_stream_conv2d_4_source_35_pat_cur_offset_3 + _source_stream_conv2d_4_source_35_pat_stride_buf_3;
        _source_stream_conv2d_4_source_35_pat_count_3 <= _source_stream_conv2d_4_source_35_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0) && (_source_stream_conv2d_4_source_35_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_35_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_35_pat_count_3 <= _source_stream_conv2d_4_source_35_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_source_ram_renable <= 0;
        _stream_conv2d_4_source_35_idle <= 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_source_ram_renable <= 0;
        _stream_conv2d_4_source_35_idle <= 1;
      end 
      if(_set_flag_507) begin
        _stream_conv2d_4_source_36_source_mode <= 5'b10;
        _stream_conv2d_4_source_36_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_507) begin
        _source_stream_conv2d_4_source_36_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_36_pat_stride_0 <= 1;
      end 
      if(_set_flag_507) begin
        _source_stream_conv2d_4_source_36_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_36_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_507) begin
        _source_stream_conv2d_4_source_36_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_36_pat_stride_2 <= 0;
      end 
      if(_set_flag_507) begin
        _source_stream_conv2d_4_source_36_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_36_pat_stride_3 <= 0;
      end 
      if(_set_flag_507) begin
        _stream_conv2d_4_source_36_source_sel <= 19;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_source_offset_buf <= _stream_conv2d_4_source_36_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_count_0 <= _source_stream_conv2d_4_source_36_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_count_1 <= _source_stream_conv2d_4_source_36_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_count_2 <= _source_stream_conv2d_4_source_36_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_count_3 <= _source_stream_conv2d_4_source_36_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_size_buf_0 <= _source_stream_conv2d_4_source_36_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_size_buf_1 <= _source_stream_conv2d_4_source_36_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_size_buf_2 <= _source_stream_conv2d_4_source_36_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_size_buf_3 <= _source_stream_conv2d_4_source_36_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_stride_buf_0 <= _source_stream_conv2d_4_source_36_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_stride_buf_1 <= _source_stream_conv2d_4_source_36_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_stride_buf_2 <= _source_stream_conv2d_4_source_36_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_stride_buf_3 <= _source_stream_conv2d_4_source_36_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_634 <= _stream_conv2d_4_source_36_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_idle <= 0;
        _stream_conv2d_4_source_36_source_ram_raddr <= _stream_conv2d_4_source_36_source_pat_all_offset;
        _stream_conv2d_4_source_36_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_0 <= _source_stream_conv2d_4_source_36_pat_cur_offset_0 + _source_stream_conv2d_4_source_36_pat_stride_buf_0;
        _source_stream_conv2d_4_source_36_pat_count_0 <= _source_stream_conv2d_4_source_36_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_4_source_36_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_36_pat_count_0 <= _source_stream_conv2d_4_source_36_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_4_source_36_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_1 <= _source_stream_conv2d_4_source_36_pat_cur_offset_1 + _source_stream_conv2d_4_source_36_pat_stride_buf_1;
        _source_stream_conv2d_4_source_36_pat_count_1 <= _source_stream_conv2d_4_source_36_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_36_pat_count_1 <= _source_stream_conv2d_4_source_36_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_2 <= _source_stream_conv2d_4_source_36_pat_cur_offset_2 + _source_stream_conv2d_4_source_36_pat_stride_buf_2;
        _source_stream_conv2d_4_source_36_pat_count_2 <= _source_stream_conv2d_4_source_36_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_36_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_36_pat_count_2 <= _source_stream_conv2d_4_source_36_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0) && (_source_stream_conv2d_4_source_36_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_3 <= _source_stream_conv2d_4_source_36_pat_cur_offset_3 + _source_stream_conv2d_4_source_36_pat_stride_buf_3;
        _source_stream_conv2d_4_source_36_pat_count_3 <= _source_stream_conv2d_4_source_36_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0) && (_source_stream_conv2d_4_source_36_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_36_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_36_pat_count_3 <= _source_stream_conv2d_4_source_36_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_source_ram_renable <= 0;
        _stream_conv2d_4_source_36_idle <= 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_source_ram_renable <= 0;
        _stream_conv2d_4_source_36_idle <= 1;
      end 
      if(_set_flag_516) begin
        _stream_conv2d_4_source_37_source_mode <= 5'b10;
        _stream_conv2d_4_source_37_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_516) begin
        _source_stream_conv2d_4_source_37_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_37_pat_stride_0 <= 1;
      end 
      if(_set_flag_516) begin
        _source_stream_conv2d_4_source_37_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_37_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_516) begin
        _source_stream_conv2d_4_source_37_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_37_pat_stride_2 <= 0;
      end 
      if(_set_flag_516) begin
        _source_stream_conv2d_4_source_37_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_37_pat_stride_3 <= 0;
      end 
      if(_set_flag_516) begin
        _stream_conv2d_4_source_37_source_sel <= 20;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_source_offset_buf <= _stream_conv2d_4_source_37_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_count_0 <= _source_stream_conv2d_4_source_37_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_count_1 <= _source_stream_conv2d_4_source_37_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_count_2 <= _source_stream_conv2d_4_source_37_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_count_3 <= _source_stream_conv2d_4_source_37_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_size_buf_0 <= _source_stream_conv2d_4_source_37_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_size_buf_1 <= _source_stream_conv2d_4_source_37_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_size_buf_2 <= _source_stream_conv2d_4_source_37_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_size_buf_3 <= _source_stream_conv2d_4_source_37_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_stride_buf_0 <= _source_stream_conv2d_4_source_37_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_stride_buf_1 <= _source_stream_conv2d_4_source_37_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_stride_buf_2 <= _source_stream_conv2d_4_source_37_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_stride_buf_3 <= _source_stream_conv2d_4_source_37_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_635 <= _stream_conv2d_4_source_37_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_idle <= 0;
        _stream_conv2d_4_source_37_source_ram_raddr <= _stream_conv2d_4_source_37_source_pat_all_offset;
        _stream_conv2d_4_source_37_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_0 <= _source_stream_conv2d_4_source_37_pat_cur_offset_0 + _source_stream_conv2d_4_source_37_pat_stride_buf_0;
        _source_stream_conv2d_4_source_37_pat_count_0 <= _source_stream_conv2d_4_source_37_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_4_source_37_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_37_pat_count_0 <= _source_stream_conv2d_4_source_37_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_4_source_37_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_1 <= _source_stream_conv2d_4_source_37_pat_cur_offset_1 + _source_stream_conv2d_4_source_37_pat_stride_buf_1;
        _source_stream_conv2d_4_source_37_pat_count_1 <= _source_stream_conv2d_4_source_37_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_37_pat_count_1 <= _source_stream_conv2d_4_source_37_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_2 <= _source_stream_conv2d_4_source_37_pat_cur_offset_2 + _source_stream_conv2d_4_source_37_pat_stride_buf_2;
        _source_stream_conv2d_4_source_37_pat_count_2 <= _source_stream_conv2d_4_source_37_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_37_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_37_pat_count_2 <= _source_stream_conv2d_4_source_37_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0) && (_source_stream_conv2d_4_source_37_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_3 <= _source_stream_conv2d_4_source_37_pat_cur_offset_3 + _source_stream_conv2d_4_source_37_pat_stride_buf_3;
        _source_stream_conv2d_4_source_37_pat_count_3 <= _source_stream_conv2d_4_source_37_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0) && (_source_stream_conv2d_4_source_37_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_37_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_37_pat_count_3 <= _source_stream_conv2d_4_source_37_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_source_ram_renable <= 0;
        _stream_conv2d_4_source_37_idle <= 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_source_ram_renable <= 0;
        _stream_conv2d_4_source_37_idle <= 1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_526 <= _set_flag_525;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_527 <= _tmp_526;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_528 <= _tmp_527;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_529 <= _tmp_528;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_530 <= _tmp_529;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_531 <= _tmp_530;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_532 <= _tmp_531;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_533 <= _tmp_532;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_534 <= _tmp_533;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_535 <= _tmp_534;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_536 <= _tmp_535;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_537 <= _tmp_536;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_538 <= _tmp_537;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_539 <= _tmp_538;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_540 <= _tmp_539;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_541 <= _tmp_540;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_542 <= _tmp_541;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_543 <= _tmp_542;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_544 <= _tmp_543;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_545 <= _tmp_544;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_546 <= _tmp_545;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_547 <= _tmp_546;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_548 <= _tmp_547;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_549 <= _tmp_548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_550 <= _tmp_549;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_551 <= _tmp_550;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_552 <= _tmp_551;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_553 <= _tmp_552;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_554 <= _tmp_553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_555 <= _tmp_554;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_556 <= _tmp_555;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_557 <= _tmp_556;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_558 <= _tmp_557;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_561 <= _tmp_560;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_562 <= _tmp_561;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_563 <= _tmp_562;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_564 <= _tmp_563;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_565 <= _tmp_564;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_566 <= _tmp_565;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_567 <= _tmp_566;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_568 <= _tmp_567;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_569 <= _tmp_568;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_570 <= _tmp_569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_571 <= _tmp_570;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_572 <= _tmp_571;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_573 <= _tmp_572;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_574 <= _tmp_573;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_575 <= _tmp_574;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_576 <= _tmp_575;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_577 <= _tmp_576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_578 <= _tmp_577;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_579 <= _tmp_578;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_580 <= _tmp_579;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_581 <= _tmp_580;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_582 <= _tmp_581;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_583 <= _tmp_582;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_584 <= _tmp_583;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_585 <= _tmp_584;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_586 <= _tmp_585;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_587 <= _tmp_586;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_588 <= _tmp_587;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_589 <= _tmp_588;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_590 <= _tmp_589;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_591 <= _tmp_590;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_592 <= _tmp_591;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_593 <= _tmp_592;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_594 <= conv2d_4_next_stream_num_ops;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_595 <= _tmp_594;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_596 <= _tmp_595;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_597 <= _tmp_596;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_598 <= _tmp_597;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_599 <= _tmp_598;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_600 <= _tmp_599;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_601 <= _tmp_600;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_602 <= _tmp_601;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_603 <= _tmp_602;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_604 <= _tmp_603;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_605 <= _tmp_604;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_606 <= _tmp_605;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_607 <= _tmp_606;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_608 <= _tmp_607;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_609 <= _tmp_608;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_610 <= _tmp_609;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_611 <= _tmp_610;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_612 <= _tmp_611;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_613 <= _tmp_612;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_614 <= _tmp_613;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_615 <= _tmp_614;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_616 <= _tmp_615;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_617 <= _tmp_616;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_618 <= _tmp_617;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_619 <= _tmp_618;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_620 <= _tmp_619;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_621 <= _tmp_620;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_622 <= _tmp_621;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_623 <= _tmp_622;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_624 <= _tmp_623;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_625 <= _tmp_624;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_626 <= _tmp_625;
      end 
      if(_tmp_558) begin
        _stream_conv2d_4_sink_50_sink_mode <= 5'b1;
        _stream_conv2d_4_sink_50_sink_offset <= _tmp_593;
        _stream_conv2d_4_sink_50_sink_size <= _tmp_626;
        _stream_conv2d_4_sink_50_sink_stride <= 1;
      end 
      if(_tmp_558) begin
        _stream_conv2d_4_sink_50_sink_sel <= 21;
      end 
      if(_stream_conv2d_4_sink_start && _stream_conv2d_4_sink_50_sink_mode & 5'b1 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_50_sink_offset_buf <= _stream_conv2d_4_sink_50_sink_offset;
        _stream_conv2d_4_sink_50_sink_size_buf <= _stream_conv2d_4_sink_50_sink_size;
        _stream_conv2d_4_sink_50_sink_stride_buf <= _stream_conv2d_4_sink_50_sink_stride;
      end 
      if((_stream_conv2d_4_sink_50_sink_fsm_20 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_50_sink_waddr <= _stream_conv2d_4_sink_50_sink_offset_buf - _stream_conv2d_4_sink_50_sink_stride_buf;
        _stream_conv2d_4_sink_50_sink_count <= _stream_conv2d_4_sink_50_sink_size_buf;
      end 
      if((_stream_conv2d_4_sink_50_sink_fsm_20 == 2) && stream_conv2d_4_sink_51_data && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_50_sink_waddr <= _stream_conv2d_4_sink_50_sink_waddr + _stream_conv2d_4_sink_50_sink_stride_buf;
        _stream_conv2d_4_sink_50_sink_wdata <= stream_conv2d_4_sink_50_data;
        _stream_conv2d_4_sink_50_sink_wenable <= 1;
        _stream_conv2d_4_sink_50_sink_count <= _stream_conv2d_4_sink_50_sink_count - 1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1017 <= _stream_conv2d_4_source_start;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1018 <= _tmp_1017;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1019 <= _tmp_1018;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1020 <= _stream_conv2d_4_source_start;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1021 <= _tmp_1020;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1022 <= _tmp_1021;
      end 
      if(_stream_conv2d_4_stream_oready && _tmp_1022) begin
        __variable_wdata_344 <= 1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1023 <= _stream_conv2d_4_source_start;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1024 <= _tmp_1023;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1025 <= _tmp_1024;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1026 <= _tmp_1025;
      end 
      if(_stream_conv2d_4_stream_oready && _tmp_1026) begin
        __variable_wdata_344 <= 0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1029 <= _tmp_1028;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1032 <= _tmp_1031;
      end 
      if(_stream_conv2d_4_stream_oready && _tmp_1032) begin
        __variable_wdata_344 <= 1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1033 <= _stream_conv2d_4_source_start;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1034 <= _tmp_1033;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1035 <= _tmp_1034;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1036 <= _tmp_1035;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1037 <= _tmp_1036;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1038 <= _tmp_1037;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1039 <= _tmp_1038;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1040 <= _tmp_1039;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1041 <= _tmp_1040;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1042 <= _tmp_1041;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1043 <= _tmp_1042;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1044 <= _tmp_1043;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1045 <= _tmp_1044;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1046 <= _tmp_1045;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1047 <= _tmp_1046;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1048 <= _tmp_1047;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1049 <= _tmp_1048;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1050 <= _tmp_1049;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1051 <= _tmp_1050;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1052 <= _tmp_1051;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1053 <= _tmp_1052;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1054 <= _tmp_1053;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1055 <= _tmp_1054;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1056 <= _tmp_1055;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1057 <= _tmp_1056;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1058 <= _tmp_1057;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1059 <= _tmp_1058;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1060 <= _tmp_1059;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1061 <= _tmp_1060;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1062 <= _tmp_1061;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1063 <= _tmp_1062;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1064 <= _tmp_1063;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1065 <= _tmp_1064;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1066 <= _stream_conv2d_4_source_stop;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1067 <= _tmp_1066;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1068 <= _tmp_1067;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1069 <= _tmp_1068;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1070 <= _tmp_1069;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1071 <= _tmp_1070;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1072 <= _tmp_1071;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1073 <= _tmp_1072;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1074 <= _tmp_1073;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1075 <= _tmp_1074;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1076 <= _tmp_1075;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1077 <= _tmp_1076;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1078 <= _tmp_1077;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1079 <= _tmp_1078;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1080 <= _tmp_1079;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1081 <= _tmp_1080;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1082 <= _tmp_1081;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1083 <= _tmp_1082;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1084 <= _tmp_1083;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1085 <= _tmp_1084;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1086 <= _tmp_1085;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1087 <= _tmp_1086;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1088 <= _tmp_1087;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1089 <= _tmp_1088;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1090 <= _tmp_1089;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1091 <= _tmp_1090;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1092 <= _tmp_1091;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1093 <= _tmp_1092;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1094 <= _tmp_1093;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1095 <= _tmp_1094;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1096 <= _tmp_1095;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1097 <= _tmp_1096;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1098 <= _tmp_1097;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1099 <= _stream_conv2d_4_source_busy;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1100 <= _tmp_1099;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1101 <= _tmp_1100;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1102 <= _tmp_1101;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1103 <= _tmp_1102;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1104 <= _tmp_1103;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1105 <= _tmp_1104;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1106 <= _tmp_1105;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1107 <= _tmp_1106;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1108 <= _tmp_1107;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1109 <= _tmp_1108;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1110 <= _tmp_1109;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1111 <= _tmp_1110;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1112 <= _tmp_1111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1113 <= _tmp_1112;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1114 <= _tmp_1113;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1115 <= _tmp_1114;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1116 <= _tmp_1115;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1117 <= _tmp_1116;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1118 <= _tmp_1117;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1119 <= _tmp_1118;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1120 <= _tmp_1119;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1121 <= _tmp_1120;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1122 <= _tmp_1121;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1123 <= _tmp_1122;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1124 <= _tmp_1123;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1125 <= _tmp_1124;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1126 <= _tmp_1125;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1127 <= _tmp_1126;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1128 <= _tmp_1127;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1129 <= _tmp_1128;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1130 <= _tmp_1129;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1131 <= _tmp_1130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1132 <= _stream_conv2d_4_sink_busy;
      end 
      if(!_stream_conv2d_4_sink_busy && _tmp_1132) begin
        _stream_conv2d_4_busy_reg <= 0;
      end 
      if(_stream_conv2d_4_source_busy) begin
        _stream_conv2d_4_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_conv2d_4_fsm_1 = 1;
  localparam _stream_conv2d_4_fsm_2 = 2;
  localparam _stream_conv2d_4_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_init;
      _stream_conv2d_4_source_start <= 0;
      _stream_conv2d_4_source_busy <= 0;
      _stream_conv2d_4_stream_ivalid <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _tmp_1019) begin
        _stream_conv2d_4_stream_ivalid <= 1;
      end 
      if(_stream_conv2d_4_stream_oready && _tmp_1029) begin
        _stream_conv2d_4_stream_ivalid <= 0;
      end 
      case(_stream_conv2d_4_fsm)
        _stream_conv2d_4_fsm_init: begin
          if(_stream_conv2d_4_run_flag) begin
            _stream_conv2d_4_source_start <= 1;
          end 
          if(_stream_conv2d_4_run_flag) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_1;
          end 
        end
        _stream_conv2d_4_fsm_1: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_start <= 0;
            _stream_conv2d_4_source_busy <= 1;
          end 
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_2;
          end 
        end
        _stream_conv2d_4_fsm_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_3;
          end 
        end
        _stream_conv2d_4_fsm_3: begin
          if(_stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3))) begin
            _stream_conv2d_4_source_busy <= 0;
          end 
          if(_stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3)) && _stream_conv2d_4_run_flag) begin
            _stream_conv2d_4_source_start <= 1;
          end 
          if(_stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3))) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_init;
          end 
          if(_stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3)) && _stream_conv2d_4_run_flag) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_6_source_1_source_ram_renable <= 0;
      _stream_max_pool_serial_6_source_1_source_fifo_deq <= 0;
      _stream_max_pool_serial_6_source_1_idle <= 1;
      _stream_max_pool_serial_6_sink_6_sink_wenable <= 0;
      _stream_max_pool_serial_6_sink_6_sink_fifo_enq <= 0;
      _stream_max_pool_serial_6_sink_7_sink_wenable <= 0;
      _stream_max_pool_serial_6_sink_7_sink_fifo_enq <= 0;
      __stream_max_pool_serial_6_stream_ivalid_1 <= 0;
      __stream_max_pool_serial_6_stream_ivalid_2 <= 0;
      __stream_max_pool_serial_6_stream_ivalid_3 <= 0;
      __stream_max_pool_serial_6_stream_ivalid_4 <= 0;
      __stream_max_pool_serial_6_stream_ivalid_5 <= 0;
      _counter_data_932 <= 1'sd0;
      _counter_count_932 <= 1'sd0;
      __delay_data_1390__variable_930 <= 0;
      __delay_data_1391_reinterpretcast_939 <= 0;
      __delay_data_1393__variable_931 <= 0;
      __delay_data_1396__variable_928 <= 0;
      __delay_data_1399_reinterpretcast_943 <= 0;
      _pointer_data_935 <= 0;
      __delay_data_1392__delay_1391_reinterpretcast_939 <= 0;
      __delay_data_1394__delay_1393__variable_931 <= 0;
      __delay_data_1397__delay_1396__variable_928 <= 0;
      __delay_data_1400__delay_1399_reinterpretcast_943 <= 0;
      _cond_data_945 <= 0;
      _cond_data_950 <= 0;
      __delay_data_1395__delay_1394__delay_1393__variable_931 <= 0;
      __delay_data_1398__delay_1397__delay_1396__variable_928 <= 0;
      _stream_max_pool_serial_6_parameter_0_next_parameter_data <= 0;
      __variable_wdata_928 <= 0;
      _stream_max_pool_serial_6_parameter_2_next_parameter_data <= 0;
      __variable_wdata_930 <= 0;
      _stream_max_pool_serial_6_source_1_source_mode <= 5'b0;
      _stream_max_pool_serial_6_source_1_source_offset <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_3 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_3 <= 0;
      _stream_max_pool_serial_6_source_1_source_sel <= 0;
      _stream_max_pool_serial_6_source_1_source_offset_buf <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_count_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_count_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_count_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_count_3 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_buf_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_buf_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_buf_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_buf_3 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_buf_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_buf_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_buf_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_buf_3 <= 0;
      __variable_wdata_929 <= 0;
      _stream_max_pool_serial_6_source_1_source_ram_raddr <= 0;
      _tmp_1194 <= 0;
      _tmp_1195 <= 0;
      _tmp_1196 <= 0;
      _tmp_1197 <= 0;
      _tmp_1198 <= 0;
      _tmp_1199 <= 0;
      _tmp_1200 <= 0;
      _tmp_1203 <= 0;
      _tmp_1204 <= 0;
      _tmp_1205 <= 0;
      _tmp_1206 <= 0;
      _tmp_1207 <= 0;
      _tmp_1208 <= 0;
      _tmp_1209 <= 0;
      _tmp_1210 <= 0;
      _tmp_1211 <= 0;
      _tmp_1212 <= 0;
      _tmp_1213 <= 0;
      _tmp_1214 <= 0;
      _tmp_1215 <= 0;
      _tmp_1216 <= 0;
      _stream_max_pool_serial_6_sink_6_sink_mode <= 5'b0;
      _stream_max_pool_serial_6_sink_6_sink_offset <= 0;
      _stream_max_pool_serial_6_sink_6_sink_size <= 0;
      _stream_max_pool_serial_6_sink_6_sink_stride <= 0;
      _stream_max_pool_serial_6_sink_6_sink_sel <= 0;
      _stream_max_pool_serial_6_sink_6_sink_offset_buf <= 0;
      _stream_max_pool_serial_6_sink_6_sink_size_buf <= 0;
      _stream_max_pool_serial_6_sink_6_sink_stride_buf <= 0;
      _stream_max_pool_serial_6_sink_6_sink_waddr <= 0;
      _stream_max_pool_serial_6_sink_6_sink_count <= 0;
      _stream_max_pool_serial_6_sink_6_sink_wdata <= 0;
      _tmp_1258 <= 0;
      _tmp_1259 <= 0;
      _tmp_1260 <= 0;
      _tmp_1261 <= 0;
      _tmp_1262 <= 0;
      _tmp_1263 <= 0;
      __variable_wdata_931 <= 0;
      _tmp_1264 <= 0;
      _tmp_1265 <= 0;
      _tmp_1266 <= 0;
      _tmp_1267 <= 0;
      _tmp_1270 <= 0;
      _tmp_1273 <= 0;
      _tmp_1274 <= 0;
      _tmp_1275 <= 0;
      _tmp_1276 <= 0;
      _tmp_1277 <= 0;
      _tmp_1278 <= 0;
      _tmp_1279 <= 0;
      _tmp_1280 <= 0;
      _tmp_1281 <= 0;
      _tmp_1282 <= 0;
      _tmp_1283 <= 0;
      _tmp_1284 <= 0;
      _tmp_1285 <= 0;
      _tmp_1286 <= 0;
      _tmp_1287 <= 0;
      _tmp_1288 <= 0;
      _tmp_1289 <= 0;
      _tmp_1290 <= 0;
      _tmp_1291 <= 0;
      _tmp_1292 <= 0;
      _tmp_1293 <= 0;
      _tmp_1294 <= 0;
      _tmp_1295 <= 0;
      _stream_max_pool_serial_6_busy_reg <= 0;
    end else begin
      if(_stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_6_source_1_source_fifo_deq <= 0;
      end 
      _stream_max_pool_serial_6_source_1_idle <= _stream_max_pool_serial_6_source_1_idle;
      if(_stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_6_sink_wenable <= 0;
        _stream_max_pool_serial_6_sink_6_sink_fifo_enq <= 0;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_7_sink_wenable <= 0;
        _stream_max_pool_serial_6_sink_7_sink_fifo_enq <= 0;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_1 <= _stream_max_pool_serial_6_stream_ivalid;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_2 <= __stream_max_pool_serial_6_stream_ivalid_1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_3 <= __stream_max_pool_serial_6_stream_ivalid_2;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_4 <= __stream_max_pool_serial_6_stream_ivalid_3;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_5 <= __stream_max_pool_serial_6_stream_ivalid_4;
      end 
      if(_stream_max_pool_serial_6_stream_ivalid && _stream_max_pool_serial_6_stream_oready && _counter_reset_cond_932) begin
        _counter_data_932 <= 1'sd0;
      end 
      if(_stream_max_pool_serial_6_stream_ivalid && _stream_max_pool_serial_6_stream_oready) begin
        _counter_data_932 <= _counter_current_count_932;
      end 
      if(_stream_max_pool_serial_6_stream_ivalid && _stream_max_pool_serial_6_stream_oready) begin
        _counter_count_932 <= (_counter_current_count_932 >= stream_max_pool_serial_6_parameter_0_data - 2'sd1)? _counter_current_count_932 + 2'sd1 - stream_max_pool_serial_6_parameter_0_data : _counter_current_count_932 + 2'sd1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_1390__variable_930 <= stream_max_pool_serial_6_parameter_2_data;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_1391_reinterpretcast_939 <= _reinterpretcast_data_939;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_1393__variable_931 <= stream_max_pool_serial_6__reduce_reset_data;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_1396__variable_928 <= stream_max_pool_serial_6_parameter_0_data;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_1399_reinterpretcast_943 <= _reinterpretcast_data_943;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _pointer_data_935 <= __delay_data_1390__variable_930[_counter_data_932];
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_1392__delay_1391_reinterpretcast_939 <= __delay_data_1391_reinterpretcast_939;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_1394__delay_1393__variable_931 <= __delay_data_1393__variable_931;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_1397__delay_1396__variable_928 <= __delay_data_1396__variable_928;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_1400__delay_1399_reinterpretcast_943 <= __delay_data_1399_reinterpretcast_943;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _cond_data_945 <= (_pointer_data_935)? -17'sd32768 : __delay_data_1392__delay_1391_reinterpretcast_939;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _cond_data_950 <= (_pointer_data_935)? -17'sd32768 : __delay_data_1400__delay_1399_reinterpretcast_943;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_1395__delay_1394__delay_1393__variable_931 <= __delay_data_1394__delay_1393__variable_931;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_1398__delay_1397__delay_1396__variable_928 <= __delay_data_1397__delay_1396__variable_928;
      end 
      if(_set_flag_1188) begin
        _stream_max_pool_serial_6_parameter_0_next_parameter_data <= 4;
      end 
      if(_stream_max_pool_serial_6_source_start) begin
        __variable_wdata_928 <= _stream_max_pool_serial_6_parameter_0_next_parameter_data;
      end 
      if(_set_flag_1189) begin
        _stream_max_pool_serial_6_parameter_2_next_parameter_data <= max_pool_serial_6_stream_pad_masks;
      end 
      if(_stream_max_pool_serial_6_source_start) begin
        __variable_wdata_930 <= _stream_max_pool_serial_6_parameter_2_next_parameter_data;
      end 
      if(_set_flag_1190) begin
        _stream_max_pool_serial_6_source_1_source_mode <= 5'b10;
        _stream_max_pool_serial_6_source_1_source_offset <= max_pool_serial_6_stream_act_local + max_pool_serial_6_act_page_comp_offset_buf;
      end 
      if(_set_flag_1190) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_0 <= 2;
        _source_stream_max_pool_serial_6_source_1_pat_stride_0 <= cparam_max_pool_serial_6_act_read_block;
      end 
      if(_set_flag_1190) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_1 <= 2;
        _source_stream_max_pool_serial_6_source_1_pat_stride_1 <= cparam_max_pool_serial_6_act_read_size;
      end 
      if(_set_flag_1190) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_2 <= cparam_max_pool_serial_6_stream_size;
        _source_stream_max_pool_serial_6_source_1_pat_stride_2 <= 1;
      end 
      if(_set_flag_1190) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_3 <= 1;
        _source_stream_max_pool_serial_6_source_1_pat_stride_3 <= 0;
      end 
      if(_set_flag_1190) begin
        _stream_max_pool_serial_6_source_1_source_sel <= 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_source_offset_buf <= _stream_max_pool_serial_6_source_1_source_offset;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 <= 0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 <= 0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 <= 0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 <= 0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_count_0 <= _source_stream_max_pool_serial_6_source_1_pat_size_0 - 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_count_1 <= _source_stream_max_pool_serial_6_source_1_pat_size_1 - 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_count_2 <= _source_stream_max_pool_serial_6_source_1_pat_size_2 - 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_count_3 <= _source_stream_max_pool_serial_6_source_1_pat_size_3 - 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_buf_0 <= _source_stream_max_pool_serial_6_source_1_pat_size_0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_buf_1 <= _source_stream_max_pool_serial_6_source_1_pat_size_1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_buf_2 <= _source_stream_max_pool_serial_6_source_1_pat_size_2;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_buf_3 <= _source_stream_max_pool_serial_6_source_1_pat_size_3;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_stride_buf_0 <= _source_stream_max_pool_serial_6_source_1_pat_stride_0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_stride_buf_1 <= _source_stream_max_pool_serial_6_source_1_pat_stride_1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_stride_buf_2 <= _source_stream_max_pool_serial_6_source_1_pat_stride_2;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_stride_buf_3 <= _source_stream_max_pool_serial_6_source_1_pat_stride_3;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_busy && _stream_max_pool_serial_6_is_root) begin
        __variable_wdata_929 <= _stream_max_pool_serial_6_source_1_source_ram_rdata;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_idle <= 0;
        _stream_max_pool_serial_6_source_1_source_ram_raddr <= _stream_max_pool_serial_6_source_1_source_pat_all_offset;
        _stream_max_pool_serial_6_source_1_source_ram_renable <= 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 <= _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 + _source_stream_max_pool_serial_6_source_1_pat_stride_buf_0;
        _source_stream_max_pool_serial_6_source_1_pat_count_0 <= _source_stream_max_pool_serial_6_source_1_pat_count_0 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 <= 0;
        _source_stream_max_pool_serial_6_source_1_pat_count_0 <= _source_stream_max_pool_serial_6_source_1_pat_size_buf_0 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 <= _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 + _source_stream_max_pool_serial_6_source_1_pat_stride_buf_1;
        _source_stream_max_pool_serial_6_source_1_pat_count_1 <= _source_stream_max_pool_serial_6_source_1_pat_count_1 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 <= 0;
        _source_stream_max_pool_serial_6_source_1_pat_count_1 <= _source_stream_max_pool_serial_6_source_1_pat_size_buf_1 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0)) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 <= _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 + _source_stream_max_pool_serial_6_source_1_pat_stride_buf_2;
        _source_stream_max_pool_serial_6_source_1_pat_count_2 <= _source_stream_max_pool_serial_6_source_1_pat_count_2 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0)) && (_source_stream_max_pool_serial_6_source_1_pat_count_2 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 <= 0;
        _source_stream_max_pool_serial_6_source_1_pat_count_2 <= _source_stream_max_pool_serial_6_source_1_pat_size_buf_2 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_2 == 0)) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 <= _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 + _source_stream_max_pool_serial_6_source_1_pat_stride_buf_3;
        _source_stream_max_pool_serial_6_source_1_pat_count_3 <= _source_stream_max_pool_serial_6_source_1_pat_count_3 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_2 == 0)) && (_source_stream_max_pool_serial_6_source_1_pat_count_3 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 <= 0;
        _source_stream_max_pool_serial_6_source_1_pat_count_3 <= _source_stream_max_pool_serial_6_source_1_pat_size_buf_3 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_6_source_stop && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_6_source_1_idle <= 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 2) && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_6_source_1_idle <= 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1194 <= _set_flag_1193;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1195 <= _tmp_1194;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1196 <= _tmp_1195;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1197 <= _tmp_1196;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1198 <= _tmp_1197;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1199 <= _tmp_1198;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1200 <= _tmp_1199;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1203 <= _tmp_1202;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1204 <= _tmp_1203;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1205 <= _tmp_1204;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1206 <= _tmp_1205;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1207 <= _tmp_1206;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1208 <= _tmp_1207;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1209 <= _tmp_1208;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1210 <= cparam_max_pool_serial_6_stream_size;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1211 <= _tmp_1210;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1212 <= _tmp_1211;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1213 <= _tmp_1212;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1214 <= _tmp_1213;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1215 <= _tmp_1214;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1216 <= _tmp_1215;
      end 
      if(_tmp_1200) begin
        _stream_max_pool_serial_6_sink_6_sink_mode <= 5'b1;
        _stream_max_pool_serial_6_sink_6_sink_offset <= _tmp_1209;
        _stream_max_pool_serial_6_sink_6_sink_size <= _tmp_1216;
        _stream_max_pool_serial_6_sink_6_sink_stride <= 1;
      end 
      if(_tmp_1200) begin
        _stream_max_pool_serial_6_sink_6_sink_sel <= 2;
      end 
      if(_stream_max_pool_serial_6_sink_start && _stream_max_pool_serial_6_sink_6_sink_mode & 5'b1 && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_6_sink_offset_buf <= _stream_max_pool_serial_6_sink_6_sink_offset;
        _stream_max_pool_serial_6_sink_6_sink_size_buf <= _stream_max_pool_serial_6_sink_6_sink_size;
        _stream_max_pool_serial_6_sink_6_sink_stride_buf <= _stream_max_pool_serial_6_sink_6_sink_stride;
      end 
      if((_stream_max_pool_serial_6_sink_6_sink_fsm_1 == 1) && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_6_sink_waddr <= _stream_max_pool_serial_6_sink_6_sink_offset_buf - _stream_max_pool_serial_6_sink_6_sink_stride_buf;
        _stream_max_pool_serial_6_sink_6_sink_count <= _stream_max_pool_serial_6_sink_6_sink_size_buf;
      end 
      if((_stream_max_pool_serial_6_sink_6_sink_fsm_1 == 2) && stream_max_pool_serial_6_sink_7_data && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_6_sink_waddr <= _stream_max_pool_serial_6_sink_6_sink_waddr + _stream_max_pool_serial_6_sink_6_sink_stride_buf;
        _stream_max_pool_serial_6_sink_6_sink_wdata <= stream_max_pool_serial_6_sink_6_data;
        _stream_max_pool_serial_6_sink_6_sink_wenable <= 1;
        _stream_max_pool_serial_6_sink_6_sink_count <= _stream_max_pool_serial_6_sink_6_sink_count - 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1258 <= _stream_max_pool_serial_6_source_start;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1259 <= _tmp_1258;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1260 <= _tmp_1259;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1261 <= _stream_max_pool_serial_6_source_start;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1262 <= _tmp_1261;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1263 <= _tmp_1262;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _tmp_1263) begin
        __variable_wdata_931 <= 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1264 <= _stream_max_pool_serial_6_source_start;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1265 <= _tmp_1264;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1266 <= _tmp_1265;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1267 <= _tmp_1266;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _tmp_1267) begin
        __variable_wdata_931 <= 0;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1270 <= _tmp_1269;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1273 <= _tmp_1272;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _tmp_1273) begin
        __variable_wdata_931 <= 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1274 <= _stream_max_pool_serial_6_source_start;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1275 <= _tmp_1274;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1276 <= _tmp_1275;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1277 <= _tmp_1276;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1278 <= _tmp_1277;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1279 <= _tmp_1278;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1280 <= _tmp_1279;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1281 <= _stream_max_pool_serial_6_source_stop;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1282 <= _tmp_1281;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1283 <= _tmp_1282;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1284 <= _tmp_1283;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1285 <= _tmp_1284;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1286 <= _tmp_1285;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1287 <= _tmp_1286;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1288 <= _stream_max_pool_serial_6_source_busy;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1289 <= _tmp_1288;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1290 <= _tmp_1289;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1291 <= _tmp_1290;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1292 <= _tmp_1291;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1293 <= _tmp_1292;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1294 <= _tmp_1293;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1295 <= _stream_max_pool_serial_6_sink_busy;
      end 
      if(!_stream_max_pool_serial_6_sink_busy && _tmp_1295) begin
        _stream_max_pool_serial_6_busy_reg <= 0;
      end 
      if(_stream_max_pool_serial_6_source_busy) begin
        _stream_max_pool_serial_6_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_max_pool_serial_6_fsm_1 = 1;
  localparam _stream_max_pool_serial_6_fsm_2 = 2;
  localparam _stream_max_pool_serial_6_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_init;
      _stream_max_pool_serial_6_source_start <= 0;
      _stream_max_pool_serial_6_source_busy <= 0;
      _stream_max_pool_serial_6_stream_ivalid <= 0;
    end else begin
      if(_stream_max_pool_serial_6_stream_oready && _tmp_1260) begin
        _stream_max_pool_serial_6_stream_ivalid <= 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _tmp_1270) begin
        _stream_max_pool_serial_6_stream_ivalid <= 0;
      end 
      case(_stream_max_pool_serial_6_fsm)
        _stream_max_pool_serial_6_fsm_init: begin
          if(_stream_max_pool_serial_6_run_flag) begin
            _stream_max_pool_serial_6_source_start <= 1;
          end 
          if(_stream_max_pool_serial_6_run_flag) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_1;
          end 
        end
        _stream_max_pool_serial_6_fsm_1: begin
          if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_start <= 0;
            _stream_max_pool_serial_6_source_busy <= 1;
          end 
          if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_2;
          end 
        end
        _stream_max_pool_serial_6_fsm_2: begin
          if(_stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_3;
          end 
        end
        _stream_max_pool_serial_6_fsm_3: begin
          if(_stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3))) begin
            _stream_max_pool_serial_6_source_busy <= 0;
          end 
          if(_stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3)) && _stream_max_pool_serial_6_run_flag) begin
            _stream_max_pool_serial_6_source_start <= 1;
          end 
          if(_stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3))) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_init;
          end 
          if(_stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3)) && _stream_max_pool_serial_6_run_flag) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_23_source_7_source_ram_renable <= 0;
      _stream_matmul_23_source_7_source_fifo_deq <= 0;
      _stream_matmul_23_source_7_idle <= 1;
      _stream_matmul_23_source_9_source_ram_renable <= 0;
      _stream_matmul_23_source_9_source_fifo_deq <= 0;
      _stream_matmul_23_source_9_idle <= 1;
      _stream_matmul_23_source_11_source_ram_renable <= 0;
      _stream_matmul_23_source_11_source_fifo_deq <= 0;
      _stream_matmul_23_source_11_idle <= 1;
      _stream_matmul_23_source_13_source_ram_renable <= 0;
      _stream_matmul_23_source_13_source_fifo_deq <= 0;
      _stream_matmul_23_source_13_idle <= 1;
      _stream_matmul_23_source_15_source_ram_renable <= 0;
      _stream_matmul_23_source_15_source_fifo_deq <= 0;
      _stream_matmul_23_source_15_idle <= 1;
      _stream_matmul_23_source_20_source_ram_renable <= 0;
      _stream_matmul_23_source_20_source_fifo_deq <= 0;
      _stream_matmul_23_source_20_idle <= 1;
      _stream_matmul_23_source_21_source_ram_renable <= 0;
      _stream_matmul_23_source_21_source_fifo_deq <= 0;
      _stream_matmul_23_source_21_idle <= 1;
      _stream_matmul_23_sink_26_sink_wenable <= 0;
      _stream_matmul_23_sink_26_sink_fifo_enq <= 0;
      _stream_matmul_23_sink_27_sink_wenable <= 0;
      _stream_matmul_23_sink_27_sink_fifo_enq <= 0;
      __stream_matmul_23_stream_ivalid_1 <= 0;
      __stream_matmul_23_stream_ivalid_2 <= 0;
      __stream_matmul_23_stream_ivalid_3 <= 0;
      __stream_matmul_23_stream_ivalid_4 <= 0;
      __stream_matmul_23_stream_ivalid_5 <= 0;
      __stream_matmul_23_stream_ivalid_6 <= 0;
      __stream_matmul_23_stream_ivalid_7 <= 0;
      __stream_matmul_23_stream_ivalid_8 <= 0;
      __stream_matmul_23_stream_ivalid_9 <= 0;
      __stream_matmul_23_stream_ivalid_10 <= 0;
      __stream_matmul_23_stream_ivalid_11 <= 0;
      __stream_matmul_23_stream_ivalid_12 <= 0;
      __stream_matmul_23_stream_ivalid_13 <= 0;
      __stream_matmul_23_stream_ivalid_14 <= 0;
      __stream_matmul_23_stream_ivalid_15 <= 0;
      __stream_matmul_23_stream_ivalid_16 <= 0;
      __stream_matmul_23_stream_ivalid_17 <= 0;
      __stream_matmul_23_stream_ivalid_18 <= 0;
      __stream_matmul_23_stream_ivalid_19 <= 0;
      __stream_matmul_23_stream_ivalid_20 <= 0;
      __stream_matmul_23_stream_ivalid_21 <= 0;
      __stream_matmul_23_stream_ivalid_22 <= 0;
      __stream_matmul_23_stream_ivalid_23 <= 0;
      __stream_matmul_23_stream_ivalid_24 <= 0;
      __stream_matmul_23_stream_ivalid_25 <= 0;
      __stream_matmul_23_stream_ivalid_26 <= 0;
      __stream_matmul_23_stream_ivalid_27 <= 0;
      __stream_matmul_23_stream_ivalid_28 <= 0;
      __stream_matmul_23_stream_ivalid_29 <= 0;
      _eq_data_1011 <= 0;
      _eq_data_1015 <= 0;
      _plus_data_1035 <= 0;
      _plus_data_1040 <= 0;
      _plus_data_1045 <= 0;
      __delay_data_1401__variable_1010 <= 0;
      __delay_data_1402_pointer_1030 <= 0;
      __delay_data_1403_reinterpretcast_1029 <= 0;
      __delay_data_1404__variable_961 <= 0;
      __delay_data_1425__variable_956 <= 0;
      __delay_data_1436_cond_977 <= 0;
      __delay_data_1453_cond_984 <= 0;
      __delay_data_1405__delay_1404__variable_961 <= 0;
      __delay_data_1415_plus_1040 <= 0;
      __delay_data_1426__delay_1425__variable_956 <= 0;
      __delay_data_1437__delay_1436_cond_977 <= 0;
      __delay_data_1454__delay_1453_cond_984 <= 0;
      __delay_data_1471_plus_1045 <= 0;
      __delay_data_1406__delay_1405__delay_1404__variable_961 <= 0;
      __delay_data_1416__delay_1415_plus_1040 <= 0;
      __delay_data_1427__delay_1426__delay_1425__variable_956 <= 0;
      __delay_data_1438__delay_1437__delay_1436_cond_977 <= 0;
      __delay_data_1455__delay_1454__delay_1453_cond_984 <= 0;
      __delay_data_1472__delay_1471_plus_1045 <= 0;
      __delay_data_1407__delay_1406__delay_1405____variable_961 <= 0;
      __delay_data_1417__delay_1416__delay_1415_plus_1040 <= 0;
      __delay_data_1428__delay_1427__delay_1426____variable_956 <= 0;
      __delay_data_1439__delay_1438__delay_1437__delay_1436_cond_977 <= 0;
      __delay_data_1456__delay_1455__delay_1454__delay_1453_cond_984 <= 0;
      __delay_data_1473__delay_1472__delay_1471_plus_1045 <= 0;
      __delay_data_1408__delay_1407__delay_1406____variable_961 <= 0;
      __delay_data_1418__delay_1417__delay_1416___plus_1040 <= 0;
      __delay_data_1429__delay_1428__delay_1427____variable_956 <= 0;
      __delay_data_1440__delay_1439__delay_1438__delay_1437___cond_977 <= 0;
      __delay_data_1457__delay_1456__delay_1455__delay_1454___cond_984 <= 0;
      __delay_data_1474__delay_1473__delay_1472___plus_1045 <= 0;
      __delay_data_1409__delay_1408__delay_1407____variable_961 <= 0;
      __delay_data_1419__delay_1418__delay_1417___plus_1040 <= 0;
      __delay_data_1430__delay_1429__delay_1428____variable_956 <= 0;
      __delay_data_1441__delay_1440__delay_1439__delay_1438___cond_977 <= 0;
      __delay_data_1458__delay_1457__delay_1456__delay_1455___cond_984 <= 0;
      __delay_data_1475__delay_1474__delay_1473___plus_1045 <= 0;
      __delay_data_1410__delay_1409__delay_1408____variable_961 <= 0;
      __delay_data_1420__delay_1419__delay_1418___plus_1040 <= 0;
      __delay_data_1431__delay_1430__delay_1429____variable_956 <= 0;
      __delay_data_1442__delay_1441__delay_1440__delay_1439___cond_977 <= 0;
      __delay_data_1459__delay_1458__delay_1457__delay_1456___cond_984 <= 0;
      __delay_data_1476__delay_1475__delay_1474___plus_1045 <= 0;
      __delay_data_1411__delay_1410__delay_1409____variable_961 <= 0;
      __delay_data_1421__delay_1420__delay_1419___plus_1040 <= 0;
      __delay_data_1432__delay_1431__delay_1430____variable_956 <= 0;
      __delay_data_1443__delay_1442__delay_1441__delay_1440___cond_977 <= 0;
      __delay_data_1460__delay_1459__delay_1458__delay_1457___cond_984 <= 0;
      __delay_data_1477__delay_1476__delay_1475___plus_1045 <= 0;
      __delay_data_1412__delay_1411__delay_1410____variable_961 <= 0;
      __delay_data_1422__delay_1421__delay_1420___plus_1040 <= 0;
      __delay_data_1433__delay_1432__delay_1431____variable_956 <= 0;
      __delay_data_1444__delay_1443__delay_1442__delay_1441___cond_977 <= 0;
      __delay_data_1461__delay_1460__delay_1459__delay_1458___cond_984 <= 0;
      __delay_data_1478__delay_1477__delay_1476___plus_1045 <= 0;
      __delay_data_1413__delay_1412__delay_1411____variable_961 <= 0;
      __delay_data_1423__delay_1422__delay_1421___plus_1040 <= 0;
      __delay_data_1434__delay_1433__delay_1432____variable_956 <= 0;
      __delay_data_1445__delay_1444__delay_1443__delay_1442___cond_977 <= 0;
      __delay_data_1462__delay_1461__delay_1460__delay_1459___cond_984 <= 0;
      __delay_data_1479__delay_1478__delay_1477___plus_1045 <= 0;
      __delay_data_1414__delay_1413__delay_1412____variable_961 <= 0;
      __delay_data_1424__delay_1423__delay_1422___plus_1040 <= 0;
      __delay_data_1435__delay_1434__delay_1433____variable_956 <= 0;
      __delay_data_1446__delay_1445__delay_1444__delay_1443___cond_977 <= 0;
      __delay_data_1463__delay_1462__delay_1461__delay_1460___cond_984 <= 0;
      __delay_data_1480__delay_1479__delay_1478___plus_1045 <= 0;
      __delay_data_1447__delay_1446__delay_1445__delay_1444___cond_977 <= 0;
      __delay_data_1464__delay_1463__delay_1462__delay_1461___cond_984 <= 0;
      __delay_data_1481__delay_1480__delay_1479___plus_1045 <= 0;
      __delay_data_1448__delay_1447__delay_1446__delay_1445___cond_977 <= 0;
      __delay_data_1465__delay_1464__delay_1463__delay_1462___cond_984 <= 0;
      __delay_data_1482__delay_1481__delay_1480___plus_1045 <= 0;
      __delay_data_1449__delay_1448__delay_1447__delay_1446___cond_977 <= 0;
      __delay_data_1466__delay_1465__delay_1464__delay_1463___cond_984 <= 0;
      __delay_data_1483__delay_1482__delay_1481___plus_1045 <= 0;
      __delay_data_1450__delay_1449__delay_1448__delay_1447___cond_977 <= 0;
      __delay_data_1467__delay_1466__delay_1465__delay_1464___cond_984 <= 0;
      __delay_data_1484__delay_1483__delay_1482___plus_1045 <= 0;
      __delay_data_1451__delay_1450__delay_1449__delay_1448___cond_977 <= 0;
      __delay_data_1468__delay_1467__delay_1466__delay_1465___cond_984 <= 0;
      __delay_data_1485__delay_1484__delay_1483___plus_1045 <= 0;
      __delay_data_1452__delay_1451__delay_1450__delay_1449___cond_977 <= 0;
      __delay_data_1469__delay_1468__delay_1467__delay_1466___cond_984 <= 0;
      __delay_data_1486__delay_1485__delay_1484___plus_1045 <= 0;
      _plus_data_1043 <= 0;
      __delay_data_1470__delay_1469__delay_1468__delay_1467___cond_984 <= 0;
      __delay_data_1487__delay_1486__delay_1485___plus_1045 <= 0;
      __delay_data_1489__substreamoutput_1042 <= 0;
      __delay_data_1490__delay_1489__substreamoutput_1042 <= 0;
      __delay_data_1491__delay_1490____substreamoutput_1042 <= 0;
      __delay_data_1492__delay_1491____substreamoutput_1042 <= 0;
      __delay_data_1493__delay_1492____substreamoutput_1042 <= 0;
      __delay_data_1494__delay_1493____substreamoutput_1042 <= 0;
      __delay_data_1495__delay_1494____substreamoutput_1042 <= 0;
      __delay_data_1496__delay_1495____substreamoutput_1042 <= 0;
      __delay_data_1497__delay_1496____substreamoutput_1042 <= 0;
      __delay_data_1498__delay_1497____substreamoutput_1042 <= 0;
      _greaterthan_data_1048 <= 0;
      __delay_data_1488__substreamoutput_1046 <= 0;
      __delay_data_1499__delay_1498____substreamoutput_1042 <= 0;
      _cond_data_1050 <= 0;
      __delay_data_1500__delay_1499____substreamoutput_1042 <= 0;
      _stream_matmul_23_parameter_0_next_parameter_data <= 0;
      __variable_wdata_956 <= 0;
      _stream_matmul_23_parameter_1_next_parameter_data <= 0;
      __variable_wdata_957 <= 0;
      _stream_matmul_23_parameter_2_next_parameter_data <= 0;
      __variable_wdata_958 <= 0;
      _stream_matmul_23_parameter_3_next_parameter_data <= 0;
      __variable_wdata_959 <= 0;
      _stream_matmul_23_parameter_4_next_parameter_data <= 0;
      __variable_wdata_960 <= 0;
      _stream_matmul_23_parameter_6_next_parameter_data <= 0;
      __variable_wdata_971 <= 0;
      _stream_matmul_23_source_7_source_mode <= 5'b0;
      _stream_matmul_23_source_7_source_offset <= 0;
      _source_stream_matmul_23_source_7_pat_size_0 <= 0;
      _source_stream_matmul_23_source_7_pat_stride_0 <= 0;
      _source_stream_matmul_23_source_7_pat_size_1 <= 0;
      _source_stream_matmul_23_source_7_pat_stride_1 <= 0;
      _source_stream_matmul_23_source_7_pat_size_2 <= 0;
      _source_stream_matmul_23_source_7_pat_stride_2 <= 0;
      _source_stream_matmul_23_source_7_pat_size_3 <= 0;
      _source_stream_matmul_23_source_7_pat_stride_3 <= 0;
      _stream_matmul_23_source_7_source_sel <= 0;
      _stream_matmul_23_source_7_source_offset_buf <= 0;
      _source_stream_matmul_23_source_7_pat_cur_offset_0 <= 0;
      _source_stream_matmul_23_source_7_pat_cur_offset_1 <= 0;
      _source_stream_matmul_23_source_7_pat_cur_offset_2 <= 0;
      _source_stream_matmul_23_source_7_pat_cur_offset_3 <= 0;
      _source_stream_matmul_23_source_7_pat_count_0 <= 0;
      _source_stream_matmul_23_source_7_pat_count_1 <= 0;
      _source_stream_matmul_23_source_7_pat_count_2 <= 0;
      _source_stream_matmul_23_source_7_pat_count_3 <= 0;
      _source_stream_matmul_23_source_7_pat_size_buf_0 <= 0;
      _source_stream_matmul_23_source_7_pat_size_buf_1 <= 0;
      _source_stream_matmul_23_source_7_pat_size_buf_2 <= 0;
      _source_stream_matmul_23_source_7_pat_size_buf_3 <= 0;
      _source_stream_matmul_23_source_7_pat_stride_buf_0 <= 0;
      _source_stream_matmul_23_source_7_pat_stride_buf_1 <= 0;
      _source_stream_matmul_23_source_7_pat_stride_buf_2 <= 0;
      _source_stream_matmul_23_source_7_pat_stride_buf_3 <= 0;
      __variable_wdata_972 <= 0;
      _stream_matmul_23_source_7_source_ram_raddr <= 0;
      _stream_matmul_23_parameter_8_next_parameter_data <= 0;
      __variable_wdata_978 <= 0;
      _stream_matmul_23_source_9_source_mode <= 5'b0;
      _stream_matmul_23_source_9_source_offset <= 0;
      _source_stream_matmul_23_source_9_pat_size_0 <= 0;
      _source_stream_matmul_23_source_9_pat_stride_0 <= 0;
      _source_stream_matmul_23_source_9_pat_size_1 <= 0;
      _source_stream_matmul_23_source_9_pat_stride_1 <= 0;
      _source_stream_matmul_23_source_9_pat_size_2 <= 0;
      _source_stream_matmul_23_source_9_pat_stride_2 <= 0;
      _source_stream_matmul_23_source_9_pat_size_3 <= 0;
      _source_stream_matmul_23_source_9_pat_stride_3 <= 0;
      _stream_matmul_23_source_9_source_sel <= 0;
      _stream_matmul_23_source_9_source_offset_buf <= 0;
      _source_stream_matmul_23_source_9_pat_cur_offset_0 <= 0;
      _source_stream_matmul_23_source_9_pat_cur_offset_1 <= 0;
      _source_stream_matmul_23_source_9_pat_cur_offset_2 <= 0;
      _source_stream_matmul_23_source_9_pat_cur_offset_3 <= 0;
      _source_stream_matmul_23_source_9_pat_count_0 <= 0;
      _source_stream_matmul_23_source_9_pat_count_1 <= 0;
      _source_stream_matmul_23_source_9_pat_count_2 <= 0;
      _source_stream_matmul_23_source_9_pat_count_3 <= 0;
      _source_stream_matmul_23_source_9_pat_size_buf_0 <= 0;
      _source_stream_matmul_23_source_9_pat_size_buf_1 <= 0;
      _source_stream_matmul_23_source_9_pat_size_buf_2 <= 0;
      _source_stream_matmul_23_source_9_pat_size_buf_3 <= 0;
      _source_stream_matmul_23_source_9_pat_stride_buf_0 <= 0;
      _source_stream_matmul_23_source_9_pat_stride_buf_1 <= 0;
      _source_stream_matmul_23_source_9_pat_stride_buf_2 <= 0;
      _source_stream_matmul_23_source_9_pat_stride_buf_3 <= 0;
      __variable_wdata_979 <= 0;
      _stream_matmul_23_source_9_source_ram_raddr <= 0;
      _stream_matmul_23_parameter_10_next_parameter_data <= 0;
      __variable_wdata_985 <= 0;
      _stream_matmul_23_source_11_source_mode <= 5'b0;
      _stream_matmul_23_source_11_source_empty_data <= 0;
      __variable_wdata_986 <= 0;
      _stream_matmul_23_parameter_12_next_parameter_data <= 0;
      __variable_wdata_992 <= 0;
      _stream_matmul_23_source_13_source_mode <= 5'b0;
      _stream_matmul_23_source_13_source_empty_data <= 0;
      __variable_wdata_993 <= 0;
      _stream_matmul_23_parameter_14_next_parameter_data <= 0;
      __variable_wdata_999 <= 0;
      _stream_matmul_23_source_15_source_mode <= 5'b0;
      _stream_matmul_23_source_15_source_empty_data <= 0;
      __variable_wdata_1000 <= 0;
      _stream_matmul_23_parameter_16_next_parameter_data <= 0;
      __variable_wdata_1006 <= 0;
      _stream_matmul_23_parameter_17_next_parameter_data <= 0;
      __variable_wdata_1007 <= 0;
      _stream_matmul_23_parameter_18_next_parameter_data <= 0;
      __variable_wdata_1008 <= 0;
      _stream_matmul_23_parameter_19_next_parameter_data <= 0;
      __variable_wdata_1009 <= 0;
      _stream_matmul_23_source_20_source_mode <= 5'b0;
      _stream_matmul_23_source_20_source_offset <= 0;
      _source_stream_matmul_23_source_20_pat_size_0 <= 0;
      _source_stream_matmul_23_source_20_pat_stride_0 <= 0;
      _source_stream_matmul_23_source_20_pat_size_1 <= 0;
      _source_stream_matmul_23_source_20_pat_stride_1 <= 0;
      _source_stream_matmul_23_source_20_pat_size_2 <= 0;
      _source_stream_matmul_23_source_20_pat_stride_2 <= 0;
      _source_stream_matmul_23_source_20_pat_size_3 <= 0;
      _source_stream_matmul_23_source_20_pat_stride_3 <= 0;
      _stream_matmul_23_source_20_source_sel <= 0;
      _stream_matmul_23_source_20_source_offset_buf <= 0;
      _source_stream_matmul_23_source_20_pat_cur_offset_0 <= 0;
      _source_stream_matmul_23_source_20_pat_cur_offset_1 <= 0;
      _source_stream_matmul_23_source_20_pat_cur_offset_2 <= 0;
      _source_stream_matmul_23_source_20_pat_cur_offset_3 <= 0;
      _source_stream_matmul_23_source_20_pat_count_0 <= 0;
      _source_stream_matmul_23_source_20_pat_count_1 <= 0;
      _source_stream_matmul_23_source_20_pat_count_2 <= 0;
      _source_stream_matmul_23_source_20_pat_count_3 <= 0;
      _source_stream_matmul_23_source_20_pat_size_buf_0 <= 0;
      _source_stream_matmul_23_source_20_pat_size_buf_1 <= 0;
      _source_stream_matmul_23_source_20_pat_size_buf_2 <= 0;
      _source_stream_matmul_23_source_20_pat_size_buf_3 <= 0;
      _source_stream_matmul_23_source_20_pat_stride_buf_0 <= 0;
      _source_stream_matmul_23_source_20_pat_stride_buf_1 <= 0;
      _source_stream_matmul_23_source_20_pat_stride_buf_2 <= 0;
      _source_stream_matmul_23_source_20_pat_stride_buf_3 <= 0;
      __variable_wdata_1010 <= 0;
      _stream_matmul_23_source_20_source_ram_raddr <= 0;
      _stream_matmul_23_source_21_source_mode <= 5'b0;
      _stream_matmul_23_source_21_source_offset <= 0;
      _source_stream_matmul_23_source_21_pat_size_0 <= 0;
      _source_stream_matmul_23_source_21_pat_stride_0 <= 0;
      _source_stream_matmul_23_source_21_pat_size_1 <= 0;
      _source_stream_matmul_23_source_21_pat_stride_1 <= 0;
      _source_stream_matmul_23_source_21_pat_size_2 <= 0;
      _source_stream_matmul_23_source_21_pat_stride_2 <= 0;
      _source_stream_matmul_23_source_21_pat_size_3 <= 0;
      _source_stream_matmul_23_source_21_pat_stride_3 <= 0;
      _stream_matmul_23_source_21_source_sel <= 0;
      _stream_matmul_23_source_21_source_offset_buf <= 0;
      _source_stream_matmul_23_source_21_pat_cur_offset_0 <= 0;
      _source_stream_matmul_23_source_21_pat_cur_offset_1 <= 0;
      _source_stream_matmul_23_source_21_pat_cur_offset_2 <= 0;
      _source_stream_matmul_23_source_21_pat_cur_offset_3 <= 0;
      _source_stream_matmul_23_source_21_pat_count_0 <= 0;
      _source_stream_matmul_23_source_21_pat_count_1 <= 0;
      _source_stream_matmul_23_source_21_pat_count_2 <= 0;
      _source_stream_matmul_23_source_21_pat_count_3 <= 0;
      _source_stream_matmul_23_source_21_pat_size_buf_0 <= 0;
      _source_stream_matmul_23_source_21_pat_size_buf_1 <= 0;
      _source_stream_matmul_23_source_21_pat_size_buf_2 <= 0;
      _source_stream_matmul_23_source_21_pat_size_buf_3 <= 0;
      _source_stream_matmul_23_source_21_pat_stride_buf_0 <= 0;
      _source_stream_matmul_23_source_21_pat_stride_buf_1 <= 0;
      _source_stream_matmul_23_source_21_pat_stride_buf_2 <= 0;
      _source_stream_matmul_23_source_21_pat_stride_buf_3 <= 0;
      __variable_wdata_1024 <= 0;
      _stream_matmul_23_source_21_source_ram_raddr <= 0;
      _tmp_1412 <= 0;
      _tmp_1413 <= 0;
      _tmp_1414 <= 0;
      _tmp_1415 <= 0;
      _tmp_1416 <= 0;
      _tmp_1417 <= 0;
      _tmp_1418 <= 0;
      _tmp_1419 <= 0;
      _tmp_1420 <= 0;
      _tmp_1421 <= 0;
      _tmp_1422 <= 0;
      _tmp_1423 <= 0;
      _tmp_1424 <= 0;
      _tmp_1425 <= 0;
      _tmp_1426 <= 0;
      _tmp_1427 <= 0;
      _tmp_1428 <= 0;
      _tmp_1429 <= 0;
      _tmp_1430 <= 0;
      _tmp_1431 <= 0;
      _tmp_1432 <= 0;
      _tmp_1433 <= 0;
      _tmp_1434 <= 0;
      _tmp_1435 <= 0;
      _tmp_1436 <= 0;
      _tmp_1437 <= 0;
      _tmp_1438 <= 0;
      _tmp_1439 <= 0;
      _tmp_1440 <= 0;
      _tmp_1441 <= 0;
      _tmp_1442 <= 0;
      _tmp_1445 <= 0;
      _tmp_1446 <= 0;
      _tmp_1447 <= 0;
      _tmp_1448 <= 0;
      _tmp_1449 <= 0;
      _tmp_1450 <= 0;
      _tmp_1451 <= 0;
      _tmp_1452 <= 0;
      _tmp_1453 <= 0;
      _tmp_1454 <= 0;
      _tmp_1455 <= 0;
      _tmp_1456 <= 0;
      _tmp_1457 <= 0;
      _tmp_1458 <= 0;
      _tmp_1459 <= 0;
      _tmp_1460 <= 0;
      _tmp_1461 <= 0;
      _tmp_1462 <= 0;
      _tmp_1463 <= 0;
      _tmp_1464 <= 0;
      _tmp_1465 <= 0;
      _tmp_1466 <= 0;
      _tmp_1467 <= 0;
      _tmp_1468 <= 0;
      _tmp_1469 <= 0;
      _tmp_1470 <= 0;
      _tmp_1471 <= 0;
      _tmp_1472 <= 0;
      _tmp_1473 <= 0;
      _tmp_1474 <= 0;
      _tmp_1475 <= 0;
      _tmp_1476 <= 0;
      _tmp_1477 <= 0;
      _tmp_1478 <= 0;
      _tmp_1479 <= 0;
      _tmp_1480 <= 0;
      _tmp_1481 <= 0;
      _tmp_1482 <= 0;
      _tmp_1483 <= 0;
      _tmp_1484 <= 0;
      _tmp_1485 <= 0;
      _tmp_1486 <= 0;
      _tmp_1487 <= 0;
      _tmp_1488 <= 0;
      _tmp_1489 <= 0;
      _tmp_1490 <= 0;
      _tmp_1491 <= 0;
      _tmp_1492 <= 0;
      _tmp_1493 <= 0;
      _tmp_1494 <= 0;
      _tmp_1495 <= 0;
      _tmp_1496 <= 0;
      _tmp_1497 <= 0;
      _tmp_1498 <= 0;
      _tmp_1499 <= 0;
      _tmp_1500 <= 0;
      _tmp_1501 <= 0;
      _tmp_1502 <= 0;
      _tmp_1503 <= 0;
      _tmp_1504 <= 0;
      _tmp_1505 <= 0;
      _tmp_1506 <= 0;
      _stream_matmul_23_sink_26_sink_mode <= 5'b0;
      _stream_matmul_23_sink_26_sink_offset <= 0;
      _stream_matmul_23_sink_26_sink_size <= 0;
      _stream_matmul_23_sink_26_sink_stride <= 0;
      _stream_matmul_23_sink_26_sink_sel <= 0;
      _stream_matmul_23_sink_26_sink_offset_buf <= 0;
      _stream_matmul_23_sink_26_sink_size_buf <= 0;
      _stream_matmul_23_sink_26_sink_stride_buf <= 0;
      _stream_matmul_23_sink_26_sink_waddr <= 0;
      _stream_matmul_23_sink_26_sink_count <= 0;
      _stream_matmul_23_sink_26_sink_wdata <= 0;
      _tmp_1519 <= 0;
      _tmp_1520 <= 0;
      _tmp_1521 <= 0;
      _tmp_1522 <= 0;
      _tmp_1523 <= 0;
      _tmp_1524 <= 0;
      __variable_wdata_961 <= 0;
      _tmp_1525 <= 0;
      _tmp_1526 <= 0;
      _tmp_1527 <= 0;
      _tmp_1528 <= 0;
      _tmp_1531 <= 0;
      _tmp_1534 <= 0;
      _tmp_1535 <= 0;
      _tmp_1536 <= 0;
      _tmp_1537 <= 0;
      _tmp_1538 <= 0;
      _tmp_1539 <= 0;
      _tmp_1540 <= 0;
      _tmp_1541 <= 0;
      _tmp_1542 <= 0;
      _tmp_1543 <= 0;
      _tmp_1544 <= 0;
      _tmp_1545 <= 0;
      _tmp_1546 <= 0;
      _tmp_1547 <= 0;
      _tmp_1548 <= 0;
      _tmp_1549 <= 0;
      _tmp_1550 <= 0;
      _tmp_1551 <= 0;
      _tmp_1552 <= 0;
      _tmp_1553 <= 0;
      _tmp_1554 <= 0;
      _tmp_1555 <= 0;
      _tmp_1556 <= 0;
      _tmp_1557 <= 0;
      _tmp_1558 <= 0;
      _tmp_1559 <= 0;
      _tmp_1560 <= 0;
      _tmp_1561 <= 0;
      _tmp_1562 <= 0;
      _tmp_1563 <= 0;
      _tmp_1564 <= 0;
      _tmp_1565 <= 0;
      _tmp_1566 <= 0;
      _tmp_1567 <= 0;
      _tmp_1568 <= 0;
      _tmp_1569 <= 0;
      _tmp_1570 <= 0;
      _tmp_1571 <= 0;
      _tmp_1572 <= 0;
      _tmp_1573 <= 0;
      _tmp_1574 <= 0;
      _tmp_1575 <= 0;
      _tmp_1576 <= 0;
      _tmp_1577 <= 0;
      _tmp_1578 <= 0;
      _tmp_1579 <= 0;
      _tmp_1580 <= 0;
      _tmp_1581 <= 0;
      _tmp_1582 <= 0;
      _tmp_1583 <= 0;
      _tmp_1584 <= 0;
      _tmp_1585 <= 0;
      _tmp_1586 <= 0;
      _tmp_1587 <= 0;
      _tmp_1588 <= 0;
      _tmp_1589 <= 0;
      _tmp_1590 <= 0;
      _tmp_1591 <= 0;
      _tmp_1592 <= 0;
      _tmp_1593 <= 0;
      _tmp_1594 <= 0;
      _tmp_1595 <= 0;
      _tmp_1596 <= 0;
      _tmp_1597 <= 0;
      _tmp_1598 <= 0;
      _tmp_1599 <= 0;
      _tmp_1600 <= 0;
      _tmp_1601 <= 0;
      _tmp_1602 <= 0;
      _tmp_1603 <= 0;
      _tmp_1604 <= 0;
      _tmp_1605 <= 0;
      _tmp_1606 <= 0;
      _tmp_1607 <= 0;
      _tmp_1608 <= 0;
      _tmp_1609 <= 0;
      _tmp_1610 <= 0;
      _tmp_1611 <= 0;
      _tmp_1612 <= 0;
      _tmp_1613 <= 0;
      _tmp_1614 <= 0;
      _tmp_1615 <= 0;
      _tmp_1616 <= 0;
      _tmp_1617 <= 0;
      _tmp_1618 <= 0;
      _tmp_1619 <= 0;
      _tmp_1620 <= 0;
      _tmp_1621 <= 0;
      _tmp_1622 <= 0;
      _tmp_1623 <= 0;
      _tmp_1624 <= 0;
      _tmp_1625 <= 0;
      _tmp_1626 <= 0;
      _tmp_1627 <= 0;
      _tmp_1628 <= 0;
      _stream_matmul_23_busy_reg <= 0;
    end else begin
      if(_stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_7_source_ram_renable <= 0;
        _stream_matmul_23_source_7_source_fifo_deq <= 0;
      end 
      _stream_matmul_23_source_7_idle <= _stream_matmul_23_source_7_idle;
      if(_stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_9_source_ram_renable <= 0;
        _stream_matmul_23_source_9_source_fifo_deq <= 0;
      end 
      _stream_matmul_23_source_9_idle <= _stream_matmul_23_source_9_idle;
      if(_stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_11_source_ram_renable <= 0;
        _stream_matmul_23_source_11_source_fifo_deq <= 0;
      end 
      _stream_matmul_23_source_11_idle <= _stream_matmul_23_source_11_idle;
      if(_stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_13_source_ram_renable <= 0;
        _stream_matmul_23_source_13_source_fifo_deq <= 0;
      end 
      _stream_matmul_23_source_13_idle <= _stream_matmul_23_source_13_idle;
      if(_stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_15_source_ram_renable <= 0;
        _stream_matmul_23_source_15_source_fifo_deq <= 0;
      end 
      _stream_matmul_23_source_15_idle <= _stream_matmul_23_source_15_idle;
      if(_stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_20_source_ram_renable <= 0;
        _stream_matmul_23_source_20_source_fifo_deq <= 0;
      end 
      _stream_matmul_23_source_20_idle <= _stream_matmul_23_source_20_idle;
      if(_stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_21_source_ram_renable <= 0;
        _stream_matmul_23_source_21_source_fifo_deq <= 0;
      end 
      _stream_matmul_23_source_21_idle <= _stream_matmul_23_source_21_idle;
      if(_stream_matmul_23_stream_oready) begin
        _stream_matmul_23_sink_26_sink_wenable <= 0;
        _stream_matmul_23_sink_26_sink_fifo_enq <= 0;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _stream_matmul_23_sink_27_sink_wenable <= 0;
        _stream_matmul_23_sink_27_sink_fifo_enq <= 0;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_1 <= _stream_matmul_23_stream_ivalid;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_2 <= __stream_matmul_23_stream_ivalid_1;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_3 <= __stream_matmul_23_stream_ivalid_2;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_4 <= __stream_matmul_23_stream_ivalid_3;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_5 <= __stream_matmul_23_stream_ivalid_4;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_6 <= __stream_matmul_23_stream_ivalid_5;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_7 <= __stream_matmul_23_stream_ivalid_6;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_8 <= __stream_matmul_23_stream_ivalid_7;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_9 <= __stream_matmul_23_stream_ivalid_8;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_10 <= __stream_matmul_23_stream_ivalid_9;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_11 <= __stream_matmul_23_stream_ivalid_10;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_12 <= __stream_matmul_23_stream_ivalid_11;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_13 <= __stream_matmul_23_stream_ivalid_12;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_14 <= __stream_matmul_23_stream_ivalid_13;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_15 <= __stream_matmul_23_stream_ivalid_14;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_16 <= __stream_matmul_23_stream_ivalid_15;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_17 <= __stream_matmul_23_stream_ivalid_16;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_18 <= __stream_matmul_23_stream_ivalid_17;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_19 <= __stream_matmul_23_stream_ivalid_18;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_20 <= __stream_matmul_23_stream_ivalid_19;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_21 <= __stream_matmul_23_stream_ivalid_20;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_22 <= __stream_matmul_23_stream_ivalid_21;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_23 <= __stream_matmul_23_stream_ivalid_22;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_24 <= __stream_matmul_23_stream_ivalid_23;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_25 <= __stream_matmul_23_stream_ivalid_24;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_26 <= __stream_matmul_23_stream_ivalid_25;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_27 <= __stream_matmul_23_stream_ivalid_26;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_28 <= __stream_matmul_23_stream_ivalid_27;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __stream_matmul_23_stream_ivalid_29 <= __stream_matmul_23_stream_ivalid_28;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _eq_data_1011 <= stream_matmul_23_parameter_1_data == 1'sd0;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _eq_data_1015 <= stream_matmul_23_parameter_2_data == 1'sd0;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _plus_data_1035 <= _cond_data_991 + stream_matmul_23_parameter_16_data;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _plus_data_1040 <= _cond_data_998 + stream_matmul_23_parameter_17_data;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _plus_data_1045 <= _cond_data_1005 + stream_matmul_23_parameter_18_data;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1401__variable_1010 <= stream_matmul_23_source_20_data;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1402_pointer_1030 <= _pointer_data_1030;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1403_reinterpretcast_1029 <= _reinterpretcast_data_1029;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1404__variable_961 <= stream_matmul_23__reduce_reset_data;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1425__variable_956 <= stream_matmul_23_parameter_0_data;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1436_cond_977 <= _cond_data_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1453_cond_984 <= _cond_data_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1405__delay_1404__variable_961 <= __delay_data_1404__variable_961;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1415_plus_1040 <= _plus_data_1040;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1426__delay_1425__variable_956 <= __delay_data_1425__variable_956;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1437__delay_1436_cond_977 <= __delay_data_1436_cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1454__delay_1453_cond_984 <= __delay_data_1453_cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1471_plus_1045 <= _plus_data_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1406__delay_1405__delay_1404__variable_961 <= __delay_data_1405__delay_1404__variable_961;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1416__delay_1415_plus_1040 <= __delay_data_1415_plus_1040;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1427__delay_1426__delay_1425__variable_956 <= __delay_data_1426__delay_1425__variable_956;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1438__delay_1437__delay_1436_cond_977 <= __delay_data_1437__delay_1436_cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1455__delay_1454__delay_1453_cond_984 <= __delay_data_1454__delay_1453_cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1472__delay_1471_plus_1045 <= __delay_data_1471_plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1407__delay_1406__delay_1405____variable_961 <= __delay_data_1406__delay_1405__delay_1404__variable_961;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1417__delay_1416__delay_1415_plus_1040 <= __delay_data_1416__delay_1415_plus_1040;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1428__delay_1427__delay_1426____variable_956 <= __delay_data_1427__delay_1426__delay_1425__variable_956;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1439__delay_1438__delay_1437__delay_1436_cond_977 <= __delay_data_1438__delay_1437__delay_1436_cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1456__delay_1455__delay_1454__delay_1453_cond_984 <= __delay_data_1455__delay_1454__delay_1453_cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1473__delay_1472__delay_1471_plus_1045 <= __delay_data_1472__delay_1471_plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1408__delay_1407__delay_1406____variable_961 <= __delay_data_1407__delay_1406__delay_1405____variable_961;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1418__delay_1417__delay_1416___plus_1040 <= __delay_data_1417__delay_1416__delay_1415_plus_1040;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1429__delay_1428__delay_1427____variable_956 <= __delay_data_1428__delay_1427__delay_1426____variable_956;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1440__delay_1439__delay_1438__delay_1437___cond_977 <= __delay_data_1439__delay_1438__delay_1437__delay_1436_cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1457__delay_1456__delay_1455__delay_1454___cond_984 <= __delay_data_1456__delay_1455__delay_1454__delay_1453_cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1474__delay_1473__delay_1472___plus_1045 <= __delay_data_1473__delay_1472__delay_1471_plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1409__delay_1408__delay_1407____variable_961 <= __delay_data_1408__delay_1407__delay_1406____variable_961;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1419__delay_1418__delay_1417___plus_1040 <= __delay_data_1418__delay_1417__delay_1416___plus_1040;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1430__delay_1429__delay_1428____variable_956 <= __delay_data_1429__delay_1428__delay_1427____variable_956;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1441__delay_1440__delay_1439__delay_1438___cond_977 <= __delay_data_1440__delay_1439__delay_1438__delay_1437___cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1458__delay_1457__delay_1456__delay_1455___cond_984 <= __delay_data_1457__delay_1456__delay_1455__delay_1454___cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1475__delay_1474__delay_1473___plus_1045 <= __delay_data_1474__delay_1473__delay_1472___plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1410__delay_1409__delay_1408____variable_961 <= __delay_data_1409__delay_1408__delay_1407____variable_961;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1420__delay_1419__delay_1418___plus_1040 <= __delay_data_1419__delay_1418__delay_1417___plus_1040;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1431__delay_1430__delay_1429____variable_956 <= __delay_data_1430__delay_1429__delay_1428____variable_956;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1442__delay_1441__delay_1440__delay_1439___cond_977 <= __delay_data_1441__delay_1440__delay_1439__delay_1438___cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1459__delay_1458__delay_1457__delay_1456___cond_984 <= __delay_data_1458__delay_1457__delay_1456__delay_1455___cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1476__delay_1475__delay_1474___plus_1045 <= __delay_data_1475__delay_1474__delay_1473___plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1411__delay_1410__delay_1409____variable_961 <= __delay_data_1410__delay_1409__delay_1408____variable_961;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1421__delay_1420__delay_1419___plus_1040 <= __delay_data_1420__delay_1419__delay_1418___plus_1040;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1432__delay_1431__delay_1430____variable_956 <= __delay_data_1431__delay_1430__delay_1429____variable_956;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1443__delay_1442__delay_1441__delay_1440___cond_977 <= __delay_data_1442__delay_1441__delay_1440__delay_1439___cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1460__delay_1459__delay_1458__delay_1457___cond_984 <= __delay_data_1459__delay_1458__delay_1457__delay_1456___cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1477__delay_1476__delay_1475___plus_1045 <= __delay_data_1476__delay_1475__delay_1474___plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1412__delay_1411__delay_1410____variable_961 <= __delay_data_1411__delay_1410__delay_1409____variable_961;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1422__delay_1421__delay_1420___plus_1040 <= __delay_data_1421__delay_1420__delay_1419___plus_1040;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1433__delay_1432__delay_1431____variable_956 <= __delay_data_1432__delay_1431__delay_1430____variable_956;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1444__delay_1443__delay_1442__delay_1441___cond_977 <= __delay_data_1443__delay_1442__delay_1441__delay_1440___cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1461__delay_1460__delay_1459__delay_1458___cond_984 <= __delay_data_1460__delay_1459__delay_1458__delay_1457___cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1478__delay_1477__delay_1476___plus_1045 <= __delay_data_1477__delay_1476__delay_1475___plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1413__delay_1412__delay_1411____variable_961 <= __delay_data_1412__delay_1411__delay_1410____variable_961;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1423__delay_1422__delay_1421___plus_1040 <= __delay_data_1422__delay_1421__delay_1420___plus_1040;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1434__delay_1433__delay_1432____variable_956 <= __delay_data_1433__delay_1432__delay_1431____variable_956;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1445__delay_1444__delay_1443__delay_1442___cond_977 <= __delay_data_1444__delay_1443__delay_1442__delay_1441___cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1462__delay_1461__delay_1460__delay_1459___cond_984 <= __delay_data_1461__delay_1460__delay_1459__delay_1458___cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1479__delay_1478__delay_1477___plus_1045 <= __delay_data_1478__delay_1477__delay_1476___plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1414__delay_1413__delay_1412____variable_961 <= __delay_data_1413__delay_1412__delay_1411____variable_961;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1424__delay_1423__delay_1422___plus_1040 <= __delay_data_1423__delay_1422__delay_1421___plus_1040;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1435__delay_1434__delay_1433____variable_956 <= __delay_data_1434__delay_1433__delay_1432____variable_956;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1446__delay_1445__delay_1444__delay_1443___cond_977 <= __delay_data_1445__delay_1444__delay_1443__delay_1442___cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1463__delay_1462__delay_1461__delay_1460___cond_984 <= __delay_data_1462__delay_1461__delay_1460__delay_1459___cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1480__delay_1479__delay_1478___plus_1045 <= __delay_data_1479__delay_1478__delay_1477___plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1447__delay_1446__delay_1445__delay_1444___cond_977 <= __delay_data_1446__delay_1445__delay_1444__delay_1443___cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1464__delay_1463__delay_1462__delay_1461___cond_984 <= __delay_data_1463__delay_1462__delay_1461__delay_1460___cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1481__delay_1480__delay_1479___plus_1045 <= __delay_data_1480__delay_1479__delay_1478___plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1448__delay_1447__delay_1446__delay_1445___cond_977 <= __delay_data_1447__delay_1446__delay_1445__delay_1444___cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1465__delay_1464__delay_1463__delay_1462___cond_984 <= __delay_data_1464__delay_1463__delay_1462__delay_1461___cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1482__delay_1481__delay_1480___plus_1045 <= __delay_data_1481__delay_1480__delay_1479___plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1449__delay_1448__delay_1447__delay_1446___cond_977 <= __delay_data_1448__delay_1447__delay_1446__delay_1445___cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1466__delay_1465__delay_1464__delay_1463___cond_984 <= __delay_data_1465__delay_1464__delay_1463__delay_1462___cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1483__delay_1482__delay_1481___plus_1045 <= __delay_data_1482__delay_1481__delay_1480___plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1450__delay_1449__delay_1448__delay_1447___cond_977 <= __delay_data_1449__delay_1448__delay_1447__delay_1446___cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1467__delay_1466__delay_1465__delay_1464___cond_984 <= __delay_data_1466__delay_1465__delay_1464__delay_1463___cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1484__delay_1483__delay_1482___plus_1045 <= __delay_data_1483__delay_1482__delay_1481___plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1451__delay_1450__delay_1449__delay_1448___cond_977 <= __delay_data_1450__delay_1449__delay_1448__delay_1447___cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1468__delay_1467__delay_1466__delay_1465___cond_984 <= __delay_data_1467__delay_1466__delay_1465__delay_1464___cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1485__delay_1484__delay_1483___plus_1045 <= __delay_data_1484__delay_1483__delay_1482___plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1452__delay_1451__delay_1450__delay_1449___cond_977 <= __delay_data_1451__delay_1450__delay_1449__delay_1448___cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1469__delay_1468__delay_1467__delay_1466___cond_984 <= __delay_data_1468__delay_1467__delay_1466__delay_1465___cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1486__delay_1485__delay_1484___plus_1045 <= __delay_data_1485__delay_1484__delay_1483___plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _plus_data_1043 <= __substreamoutput_data_1041 + __delay_data_1452__delay_1451__delay_1450__delay_1449___cond_977;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1470__delay_1469__delay_1468__delay_1467___cond_984 <= __delay_data_1469__delay_1468__delay_1467__delay_1466___cond_984;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1487__delay_1486__delay_1485___plus_1045 <= __delay_data_1486__delay_1485__delay_1484___plus_1045;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1489__substreamoutput_1042 <= __substreamoutput_data_1042;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1490__delay_1489__substreamoutput_1042 <= __delay_data_1489__substreamoutput_1042;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1491__delay_1490____substreamoutput_1042 <= __delay_data_1490__delay_1489__substreamoutput_1042;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1492__delay_1491____substreamoutput_1042 <= __delay_data_1491__delay_1490____substreamoutput_1042;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1493__delay_1492____substreamoutput_1042 <= __delay_data_1492__delay_1491____substreamoutput_1042;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1494__delay_1493____substreamoutput_1042 <= __delay_data_1493__delay_1492____substreamoutput_1042;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1495__delay_1494____substreamoutput_1042 <= __delay_data_1494__delay_1493____substreamoutput_1042;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1496__delay_1495____substreamoutput_1042 <= __delay_data_1495__delay_1494____substreamoutput_1042;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1497__delay_1496____substreamoutput_1042 <= __delay_data_1496__delay_1495____substreamoutput_1042;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1498__delay_1497____substreamoutput_1042 <= __delay_data_1497__delay_1496____substreamoutput_1042;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _greaterthan_data_1048 <= __substreamoutput_data_1046 > 1'sd0;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1488__substreamoutput_1046 <= __substreamoutput_data_1046;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1499__delay_1498____substreamoutput_1042 <= __delay_data_1498__delay_1497____substreamoutput_1042;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _cond_data_1050 <= (_greaterthan_data_1048)? __delay_data_1488__substreamoutput_1046 : 1'sd0;
      end 
      if(_stream_matmul_23_stream_oready) begin
        __delay_data_1500__delay_1499____substreamoutput_1042 <= __delay_data_1499__delay_1498____substreamoutput_1042;
      end 
      if(_set_flag_1358) begin
        _stream_matmul_23_parameter_0_next_parameter_data <= cparam_matmul_23_stream_reduce_size;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_956 <= _stream_matmul_23_parameter_0_next_parameter_data;
      end 
      if(_set_flag_1359) begin
        _stream_matmul_23_parameter_1_next_parameter_data <= matmul_23_col_select;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_957 <= _stream_matmul_23_parameter_1_next_parameter_data;
      end 
      if(_set_flag_1360) begin
        _stream_matmul_23_parameter_2_next_parameter_data <= matmul_23_row_select_buf;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_958 <= _stream_matmul_23_parameter_2_next_parameter_data;
      end 
      if(_set_flag_1361) begin
        _stream_matmul_23_parameter_3_next_parameter_data <= matmul_23_stream_pad_masks;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_959 <= _stream_matmul_23_parameter_3_next_parameter_data;
      end 
      if(_set_flag_1362) begin
        _stream_matmul_23_parameter_4_next_parameter_data <= cparam_matmul_23_stream_omit_mask;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_960 <= _stream_matmul_23_parameter_4_next_parameter_data;
      end 
      if(_set_flag_1363) begin
        _stream_matmul_23_parameter_6_next_parameter_data <= cparam_matmul_23_bias_scala;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_971 <= _stream_matmul_23_parameter_6_next_parameter_data;
      end 
      if(_set_flag_1364) begin
        _stream_matmul_23_source_7_source_mode <= 5'b10;
        _stream_matmul_23_source_7_source_offset <= (cparam_matmul_23_bias_num == 1)? 0 : matmul_23_och_count_buf;
      end 
      if(_set_flag_1364) begin
        _source_stream_matmul_23_source_7_pat_size_0 <= cparam_matmul_23_stream_reduce_size;
        _source_stream_matmul_23_source_7_pat_stride_0 <= 0;
      end 
      if(_set_flag_1364) begin
        _source_stream_matmul_23_source_7_pat_size_1 <= matmul_23_next_stream_num_ops;
        _source_stream_matmul_23_source_7_pat_stride_1 <= (cparam_matmul_23_bias_num == 1)? 0 : 1;
      end 
      if(_set_flag_1364) begin
        _source_stream_matmul_23_source_7_pat_size_2 <= 1;
        _source_stream_matmul_23_source_7_pat_stride_2 <= 0;
      end 
      if(_set_flag_1364) begin
        _source_stream_matmul_23_source_7_pat_size_3 <= 1;
        _source_stream_matmul_23_source_7_pat_stride_3 <= 0;
      end 
      if(_set_flag_1364) begin
        _stream_matmul_23_source_7_source_sel <= 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_7_source_offset_buf <= _stream_matmul_23_source_7_source_offset;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_count_0 <= _source_stream_matmul_23_source_7_pat_size_0 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_count_1 <= _source_stream_matmul_23_source_7_pat_size_1 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_count_2 <= _source_stream_matmul_23_source_7_pat_size_2 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_count_3 <= _source_stream_matmul_23_source_7_pat_size_3 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_size_buf_0 <= _source_stream_matmul_23_source_7_pat_size_0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_size_buf_1 <= _source_stream_matmul_23_source_7_pat_size_1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_size_buf_2 <= _source_stream_matmul_23_source_7_pat_size_2;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_size_buf_3 <= _source_stream_matmul_23_source_7_pat_size_3;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_stride_buf_0 <= _source_stream_matmul_23_source_7_pat_stride_0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_stride_buf_1 <= _source_stream_matmul_23_source_7_pat_stride_1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_stride_buf_2 <= _source_stream_matmul_23_source_7_pat_stride_2;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_stride_buf_3 <= _source_stream_matmul_23_source_7_pat_stride_3;
      end 
      if(_stream_matmul_23_stream_oready && _stream_matmul_23_source_busy && _stream_matmul_23_is_root) begin
        __variable_wdata_972 <= _stream_matmul_23_source_7_source_ram_rdata;
      end 
      if((_stream_matmul_23_source_7_source_pat_fsm_0 == 1) && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_7_idle <= 0;
        _stream_matmul_23_source_7_source_ram_raddr <= _stream_matmul_23_source_7_source_pat_all_offset;
        _stream_matmul_23_source_7_source_ram_renable <= 1;
      end 
      if((_stream_matmul_23_source_7_source_pat_fsm_0 == 1) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_cur_offset_0 <= _source_stream_matmul_23_source_7_pat_cur_offset_0 + _source_stream_matmul_23_source_7_pat_stride_buf_0;
        _source_stream_matmul_23_source_7_pat_count_0 <= _source_stream_matmul_23_source_7_pat_count_0 - 1;
      end 
      if((_stream_matmul_23_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_23_source_7_pat_count_0 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_cur_offset_0 <= 0;
        _source_stream_matmul_23_source_7_pat_count_0 <= _source_stream_matmul_23_source_7_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_23_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_23_source_7_pat_count_0 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_cur_offset_1 <= _source_stream_matmul_23_source_7_pat_cur_offset_1 + _source_stream_matmul_23_source_7_pat_stride_buf_1;
        _source_stream_matmul_23_source_7_pat_count_1 <= _source_stream_matmul_23_source_7_pat_count_1 - 1;
      end 
      if((_stream_matmul_23_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_23_source_7_pat_count_0 == 0) && (_source_stream_matmul_23_source_7_pat_count_1 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_cur_offset_1 <= 0;
        _source_stream_matmul_23_source_7_pat_count_1 <= _source_stream_matmul_23_source_7_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_23_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_23_source_7_pat_count_0 == 0) && (_source_stream_matmul_23_source_7_pat_count_1 == 0)) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_cur_offset_2 <= _source_stream_matmul_23_source_7_pat_cur_offset_2 + _source_stream_matmul_23_source_7_pat_stride_buf_2;
        _source_stream_matmul_23_source_7_pat_count_2 <= _source_stream_matmul_23_source_7_pat_count_2 - 1;
      end 
      if((_stream_matmul_23_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_23_source_7_pat_count_0 == 0) && (_source_stream_matmul_23_source_7_pat_count_1 == 0)) && (_source_stream_matmul_23_source_7_pat_count_2 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_cur_offset_2 <= 0;
        _source_stream_matmul_23_source_7_pat_count_2 <= _source_stream_matmul_23_source_7_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_23_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_23_source_7_pat_count_0 == 0) && (_source_stream_matmul_23_source_7_pat_count_1 == 0) && (_source_stream_matmul_23_source_7_pat_count_2 == 0)) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_cur_offset_3 <= _source_stream_matmul_23_source_7_pat_cur_offset_3 + _source_stream_matmul_23_source_7_pat_stride_buf_3;
        _source_stream_matmul_23_source_7_pat_count_3 <= _source_stream_matmul_23_source_7_pat_count_3 - 1;
      end 
      if((_stream_matmul_23_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_23_source_7_pat_count_0 == 0) && (_source_stream_matmul_23_source_7_pat_count_1 == 0) && (_source_stream_matmul_23_source_7_pat_count_2 == 0)) && (_source_stream_matmul_23_source_7_pat_count_3 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_7_pat_cur_offset_3 <= 0;
        _source_stream_matmul_23_source_7_pat_count_3 <= _source_stream_matmul_23_source_7_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_23_source_7_source_pat_fsm_0 == 1) && _stream_matmul_23_source_stop && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_7_source_ram_renable <= 0;
        _stream_matmul_23_source_7_idle <= 1;
      end 
      if((_stream_matmul_23_source_7_source_pat_fsm_0 == 2) && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_7_source_ram_renable <= 0;
        _stream_matmul_23_source_7_idle <= 1;
      end 
      if(_set_flag_1373) begin
        _stream_matmul_23_parameter_8_next_parameter_data <= cparam_matmul_23_scale_scala;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_978 <= _stream_matmul_23_parameter_8_next_parameter_data;
      end 
      if(_set_flag_1374) begin
        _stream_matmul_23_source_9_source_mode <= 5'b10;
        _stream_matmul_23_source_9_source_offset <= (cparam_matmul_23_scale_num == 1)? 0 : matmul_23_och_count_buf;
      end 
      if(_set_flag_1374) begin
        _source_stream_matmul_23_source_9_pat_size_0 <= cparam_matmul_23_stream_reduce_size;
        _source_stream_matmul_23_source_9_pat_stride_0 <= 0;
      end 
      if(_set_flag_1374) begin
        _source_stream_matmul_23_source_9_pat_size_1 <= matmul_23_next_stream_num_ops;
        _source_stream_matmul_23_source_9_pat_stride_1 <= (cparam_matmul_23_scale_num == 1)? 0 : 1;
      end 
      if(_set_flag_1374) begin
        _source_stream_matmul_23_source_9_pat_size_2 <= 1;
        _source_stream_matmul_23_source_9_pat_stride_2 <= 0;
      end 
      if(_set_flag_1374) begin
        _source_stream_matmul_23_source_9_pat_size_3 <= 1;
        _source_stream_matmul_23_source_9_pat_stride_3 <= 0;
      end 
      if(_set_flag_1374) begin
        _stream_matmul_23_source_9_source_sel <= 2;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_9_source_offset_buf <= _stream_matmul_23_source_9_source_offset;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_count_0 <= _source_stream_matmul_23_source_9_pat_size_0 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_count_1 <= _source_stream_matmul_23_source_9_pat_size_1 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_count_2 <= _source_stream_matmul_23_source_9_pat_size_2 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_count_3 <= _source_stream_matmul_23_source_9_pat_size_3 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_size_buf_0 <= _source_stream_matmul_23_source_9_pat_size_0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_size_buf_1 <= _source_stream_matmul_23_source_9_pat_size_1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_size_buf_2 <= _source_stream_matmul_23_source_9_pat_size_2;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_size_buf_3 <= _source_stream_matmul_23_source_9_pat_size_3;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_stride_buf_0 <= _source_stream_matmul_23_source_9_pat_stride_0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_stride_buf_1 <= _source_stream_matmul_23_source_9_pat_stride_1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_stride_buf_2 <= _source_stream_matmul_23_source_9_pat_stride_2;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_stride_buf_3 <= _source_stream_matmul_23_source_9_pat_stride_3;
      end 
      if(_stream_matmul_23_stream_oready && _stream_matmul_23_source_busy && _stream_matmul_23_is_root) begin
        __variable_wdata_979 <= _stream_matmul_23_source_9_source_ram_rdata;
      end 
      if((_stream_matmul_23_source_9_source_pat_fsm_1 == 1) && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_9_idle <= 0;
        _stream_matmul_23_source_9_source_ram_raddr <= _stream_matmul_23_source_9_source_pat_all_offset;
        _stream_matmul_23_source_9_source_ram_renable <= 1;
      end 
      if((_stream_matmul_23_source_9_source_pat_fsm_1 == 1) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_cur_offset_0 <= _source_stream_matmul_23_source_9_pat_cur_offset_0 + _source_stream_matmul_23_source_9_pat_stride_buf_0;
        _source_stream_matmul_23_source_9_pat_count_0 <= _source_stream_matmul_23_source_9_pat_count_0 - 1;
      end 
      if((_stream_matmul_23_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_23_source_9_pat_count_0 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_cur_offset_0 <= 0;
        _source_stream_matmul_23_source_9_pat_count_0 <= _source_stream_matmul_23_source_9_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_23_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_23_source_9_pat_count_0 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_cur_offset_1 <= _source_stream_matmul_23_source_9_pat_cur_offset_1 + _source_stream_matmul_23_source_9_pat_stride_buf_1;
        _source_stream_matmul_23_source_9_pat_count_1 <= _source_stream_matmul_23_source_9_pat_count_1 - 1;
      end 
      if((_stream_matmul_23_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_23_source_9_pat_count_0 == 0) && (_source_stream_matmul_23_source_9_pat_count_1 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_cur_offset_1 <= 0;
        _source_stream_matmul_23_source_9_pat_count_1 <= _source_stream_matmul_23_source_9_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_23_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_23_source_9_pat_count_0 == 0) && (_source_stream_matmul_23_source_9_pat_count_1 == 0)) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_cur_offset_2 <= _source_stream_matmul_23_source_9_pat_cur_offset_2 + _source_stream_matmul_23_source_9_pat_stride_buf_2;
        _source_stream_matmul_23_source_9_pat_count_2 <= _source_stream_matmul_23_source_9_pat_count_2 - 1;
      end 
      if((_stream_matmul_23_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_23_source_9_pat_count_0 == 0) && (_source_stream_matmul_23_source_9_pat_count_1 == 0)) && (_source_stream_matmul_23_source_9_pat_count_2 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_cur_offset_2 <= 0;
        _source_stream_matmul_23_source_9_pat_count_2 <= _source_stream_matmul_23_source_9_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_23_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_23_source_9_pat_count_0 == 0) && (_source_stream_matmul_23_source_9_pat_count_1 == 0) && (_source_stream_matmul_23_source_9_pat_count_2 == 0)) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_cur_offset_3 <= _source_stream_matmul_23_source_9_pat_cur_offset_3 + _source_stream_matmul_23_source_9_pat_stride_buf_3;
        _source_stream_matmul_23_source_9_pat_count_3 <= _source_stream_matmul_23_source_9_pat_count_3 - 1;
      end 
      if((_stream_matmul_23_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_23_source_9_pat_count_0 == 0) && (_source_stream_matmul_23_source_9_pat_count_1 == 0) && (_source_stream_matmul_23_source_9_pat_count_2 == 0)) && (_source_stream_matmul_23_source_9_pat_count_3 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_9_pat_cur_offset_3 <= 0;
        _source_stream_matmul_23_source_9_pat_count_3 <= _source_stream_matmul_23_source_9_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_23_source_9_source_pat_fsm_1 == 1) && _stream_matmul_23_source_stop && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_9_source_ram_renable <= 0;
        _stream_matmul_23_source_9_idle <= 1;
      end 
      if((_stream_matmul_23_source_9_source_pat_fsm_1 == 2) && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_9_source_ram_renable <= 0;
        _stream_matmul_23_source_9_idle <= 1;
      end 
      if(_set_flag_1383) begin
        _stream_matmul_23_parameter_10_next_parameter_data <= 1;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_985 <= _stream_matmul_23_parameter_10_next_parameter_data;
      end 
      if(_set_flag_1384) begin
        _stream_matmul_23_source_11_source_mode <= 5'b0;
        _stream_matmul_23_source_11_source_empty_data <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_stream_oready && !(|(_stream_matmul_23_source_11_source_mode & 5'b0))) begin
        _stream_matmul_23_source_11_idle <= 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_stream_oready && !(|(_stream_matmul_23_source_11_source_mode & 5'b0)) && _stream_matmul_23_is_root) begin
        __variable_wdata_986 <= _stream_matmul_23_source_11_source_empty_data;
      end 
      if(_set_flag_1385) begin
        _stream_matmul_23_parameter_12_next_parameter_data <= 1;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_992 <= _stream_matmul_23_parameter_12_next_parameter_data;
      end 
      if(_set_flag_1386) begin
        _stream_matmul_23_source_13_source_mode <= 5'b0;
        _stream_matmul_23_source_13_source_empty_data <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_stream_oready && !(|(_stream_matmul_23_source_13_source_mode & 5'b0))) begin
        _stream_matmul_23_source_13_idle <= 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_stream_oready && !(|(_stream_matmul_23_source_13_source_mode & 5'b0)) && _stream_matmul_23_is_root) begin
        __variable_wdata_993 <= _stream_matmul_23_source_13_source_empty_data;
      end 
      if(_set_flag_1387) begin
        _stream_matmul_23_parameter_14_next_parameter_data <= 1;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_999 <= _stream_matmul_23_parameter_14_next_parameter_data;
      end 
      if(_set_flag_1388) begin
        _stream_matmul_23_source_15_source_mode <= 5'b0;
        _stream_matmul_23_source_15_source_empty_data <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_stream_oready && !(|(_stream_matmul_23_source_15_source_mode & 5'b0))) begin
        _stream_matmul_23_source_15_idle <= 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_stream_oready && !(|(_stream_matmul_23_source_15_source_mode & 5'b0)) && _stream_matmul_23_is_root) begin
        __variable_wdata_1000 <= _stream_matmul_23_source_15_source_empty_data;
      end 
      if(_set_flag_1389) begin
        _stream_matmul_23_parameter_16_next_parameter_data <= cparam_matmul_23_cshamt_mul_value;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_1006 <= _stream_matmul_23_parameter_16_next_parameter_data;
      end 
      if(_set_flag_1390) begin
        _stream_matmul_23_parameter_17_next_parameter_data <= cparam_matmul_23_cshamt_sum_value;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_1007 <= _stream_matmul_23_parameter_17_next_parameter_data;
      end 
      if(_set_flag_1391) begin
        _stream_matmul_23_parameter_18_next_parameter_data <= cparam_matmul_23_cshamt_out_value;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_1008 <= _stream_matmul_23_parameter_18_next_parameter_data;
      end 
      if(_set_flag_1392) begin
        _stream_matmul_23_parameter_19_next_parameter_data <= cparam_matmul_23_act_func_index;
      end 
      if(_stream_matmul_23_source_start) begin
        __variable_wdata_1009 <= _stream_matmul_23_parameter_19_next_parameter_data;
      end 
      if(_set_flag_1393) begin
        _stream_matmul_23_source_20_source_mode <= 5'b10;
        _stream_matmul_23_source_20_source_offset <= matmul_23_stream_act_local_0 + matmul_23_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_1393) begin
        _source_stream_matmul_23_source_20_pat_size_0 <= cparam_matmul_23_stream_reduce_size;
        _source_stream_matmul_23_source_20_pat_stride_0 <= 1;
      end 
      if(_set_flag_1393) begin
        _source_stream_matmul_23_source_20_pat_size_1 <= matmul_23_next_stream_num_ops;
        _source_stream_matmul_23_source_20_pat_stride_1 <= 0;
      end 
      if(_set_flag_1393) begin
        _source_stream_matmul_23_source_20_pat_size_2 <= 1;
        _source_stream_matmul_23_source_20_pat_stride_2 <= 0;
      end 
      if(_set_flag_1393) begin
        _source_stream_matmul_23_source_20_pat_size_3 <= 1;
        _source_stream_matmul_23_source_20_pat_stride_3 <= 0;
      end 
      if(_set_flag_1393) begin
        _stream_matmul_23_source_20_source_sel <= 3;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_20_source_offset_buf <= _stream_matmul_23_source_20_source_offset;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_count_0 <= _source_stream_matmul_23_source_20_pat_size_0 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_count_1 <= _source_stream_matmul_23_source_20_pat_size_1 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_count_2 <= _source_stream_matmul_23_source_20_pat_size_2 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_count_3 <= _source_stream_matmul_23_source_20_pat_size_3 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_size_buf_0 <= _source_stream_matmul_23_source_20_pat_size_0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_size_buf_1 <= _source_stream_matmul_23_source_20_pat_size_1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_size_buf_2 <= _source_stream_matmul_23_source_20_pat_size_2;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_size_buf_3 <= _source_stream_matmul_23_source_20_pat_size_3;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_stride_buf_0 <= _source_stream_matmul_23_source_20_pat_stride_0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_stride_buf_1 <= _source_stream_matmul_23_source_20_pat_stride_1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_stride_buf_2 <= _source_stream_matmul_23_source_20_pat_stride_2;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_stride_buf_3 <= _source_stream_matmul_23_source_20_pat_stride_3;
      end 
      if(_stream_matmul_23_stream_oready && _stream_matmul_23_source_busy && _stream_matmul_23_is_root) begin
        __variable_wdata_1010 <= _stream_matmul_23_source_20_source_ram_rdata;
      end 
      if((_stream_matmul_23_source_20_source_pat_fsm_2 == 1) && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_20_idle <= 0;
        _stream_matmul_23_source_20_source_ram_raddr <= _stream_matmul_23_source_20_source_pat_all_offset;
        _stream_matmul_23_source_20_source_ram_renable <= 1;
      end 
      if((_stream_matmul_23_source_20_source_pat_fsm_2 == 1) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_cur_offset_0 <= _source_stream_matmul_23_source_20_pat_cur_offset_0 + _source_stream_matmul_23_source_20_pat_stride_buf_0;
        _source_stream_matmul_23_source_20_pat_count_0 <= _source_stream_matmul_23_source_20_pat_count_0 - 1;
      end 
      if((_stream_matmul_23_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_23_source_20_pat_count_0 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_cur_offset_0 <= 0;
        _source_stream_matmul_23_source_20_pat_count_0 <= _source_stream_matmul_23_source_20_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_23_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_23_source_20_pat_count_0 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_cur_offset_1 <= _source_stream_matmul_23_source_20_pat_cur_offset_1 + _source_stream_matmul_23_source_20_pat_stride_buf_1;
        _source_stream_matmul_23_source_20_pat_count_1 <= _source_stream_matmul_23_source_20_pat_count_1 - 1;
      end 
      if((_stream_matmul_23_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_23_source_20_pat_count_0 == 0) && (_source_stream_matmul_23_source_20_pat_count_1 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_cur_offset_1 <= 0;
        _source_stream_matmul_23_source_20_pat_count_1 <= _source_stream_matmul_23_source_20_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_23_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_23_source_20_pat_count_0 == 0) && (_source_stream_matmul_23_source_20_pat_count_1 == 0)) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_cur_offset_2 <= _source_stream_matmul_23_source_20_pat_cur_offset_2 + _source_stream_matmul_23_source_20_pat_stride_buf_2;
        _source_stream_matmul_23_source_20_pat_count_2 <= _source_stream_matmul_23_source_20_pat_count_2 - 1;
      end 
      if((_stream_matmul_23_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_23_source_20_pat_count_0 == 0) && (_source_stream_matmul_23_source_20_pat_count_1 == 0)) && (_source_stream_matmul_23_source_20_pat_count_2 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_cur_offset_2 <= 0;
        _source_stream_matmul_23_source_20_pat_count_2 <= _source_stream_matmul_23_source_20_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_23_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_23_source_20_pat_count_0 == 0) && (_source_stream_matmul_23_source_20_pat_count_1 == 0) && (_source_stream_matmul_23_source_20_pat_count_2 == 0)) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_cur_offset_3 <= _source_stream_matmul_23_source_20_pat_cur_offset_3 + _source_stream_matmul_23_source_20_pat_stride_buf_3;
        _source_stream_matmul_23_source_20_pat_count_3 <= _source_stream_matmul_23_source_20_pat_count_3 - 1;
      end 
      if((_stream_matmul_23_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_23_source_20_pat_count_0 == 0) && (_source_stream_matmul_23_source_20_pat_count_1 == 0) && (_source_stream_matmul_23_source_20_pat_count_2 == 0)) && (_source_stream_matmul_23_source_20_pat_count_3 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_20_pat_cur_offset_3 <= 0;
        _source_stream_matmul_23_source_20_pat_count_3 <= _source_stream_matmul_23_source_20_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_23_source_20_source_pat_fsm_2 == 1) && _stream_matmul_23_source_stop && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_20_source_ram_renable <= 0;
        _stream_matmul_23_source_20_idle <= 1;
      end 
      if((_stream_matmul_23_source_20_source_pat_fsm_2 == 2) && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_20_source_ram_renable <= 0;
        _stream_matmul_23_source_20_idle <= 1;
      end 
      if(_set_flag_1402) begin
        _stream_matmul_23_source_21_source_mode <= 5'b10;
        _stream_matmul_23_source_21_source_offset <= matmul_23_filter_page_comp_offset_buf;
      end 
      if(_set_flag_1402) begin
        _source_stream_matmul_23_source_21_pat_size_0 <= cparam_matmul_23_stream_reduce_size;
        _source_stream_matmul_23_source_21_pat_stride_0 <= 1;
      end 
      if(_set_flag_1402) begin
        _source_stream_matmul_23_source_21_pat_size_1 <= matmul_23_next_stream_num_ops;
        _source_stream_matmul_23_source_21_pat_stride_1 <= cparam_matmul_23_stream_aligned_reduce_size;
      end 
      if(_set_flag_1402) begin
        _source_stream_matmul_23_source_21_pat_size_2 <= 1;
        _source_stream_matmul_23_source_21_pat_stride_2 <= 0;
      end 
      if(_set_flag_1402) begin
        _source_stream_matmul_23_source_21_pat_size_3 <= 1;
        _source_stream_matmul_23_source_21_pat_stride_3 <= 0;
      end 
      if(_set_flag_1402) begin
        _stream_matmul_23_source_21_source_sel <= 4;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_21_source_offset_buf <= _stream_matmul_23_source_21_source_offset;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_count_0 <= _source_stream_matmul_23_source_21_pat_size_0 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_count_1 <= _source_stream_matmul_23_source_21_pat_size_1 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_count_2 <= _source_stream_matmul_23_source_21_pat_size_2 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_count_3 <= _source_stream_matmul_23_source_21_pat_size_3 - 1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_size_buf_0 <= _source_stream_matmul_23_source_21_pat_size_0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_size_buf_1 <= _source_stream_matmul_23_source_21_pat_size_1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_size_buf_2 <= _source_stream_matmul_23_source_21_pat_size_2;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_size_buf_3 <= _source_stream_matmul_23_source_21_pat_size_3;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_stride_buf_0 <= _source_stream_matmul_23_source_21_pat_stride_0;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_stride_buf_1 <= _source_stream_matmul_23_source_21_pat_stride_1;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_stride_buf_2 <= _source_stream_matmul_23_source_21_pat_stride_2;
      end 
      if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_stride_buf_3 <= _source_stream_matmul_23_source_21_pat_stride_3;
      end 
      if(_stream_matmul_23_stream_oready && _stream_matmul_23_source_busy && _stream_matmul_23_is_root) begin
        __variable_wdata_1024 <= _stream_matmul_23_source_21_source_ram_rdata;
      end 
      if((_stream_matmul_23_source_21_source_pat_fsm_3 == 1) && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_21_idle <= 0;
        _stream_matmul_23_source_21_source_ram_raddr <= _stream_matmul_23_source_21_source_pat_all_offset;
        _stream_matmul_23_source_21_source_ram_renable <= 1;
      end 
      if((_stream_matmul_23_source_21_source_pat_fsm_3 == 1) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_cur_offset_0 <= _source_stream_matmul_23_source_21_pat_cur_offset_0 + _source_stream_matmul_23_source_21_pat_stride_buf_0;
        _source_stream_matmul_23_source_21_pat_count_0 <= _source_stream_matmul_23_source_21_pat_count_0 - 1;
      end 
      if((_stream_matmul_23_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_23_source_21_pat_count_0 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_cur_offset_0 <= 0;
        _source_stream_matmul_23_source_21_pat_count_0 <= _source_stream_matmul_23_source_21_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_23_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_23_source_21_pat_count_0 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_cur_offset_1 <= _source_stream_matmul_23_source_21_pat_cur_offset_1 + _source_stream_matmul_23_source_21_pat_stride_buf_1;
        _source_stream_matmul_23_source_21_pat_count_1 <= _source_stream_matmul_23_source_21_pat_count_1 - 1;
      end 
      if((_stream_matmul_23_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_23_source_21_pat_count_0 == 0) && (_source_stream_matmul_23_source_21_pat_count_1 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_cur_offset_1 <= 0;
        _source_stream_matmul_23_source_21_pat_count_1 <= _source_stream_matmul_23_source_21_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_23_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_23_source_21_pat_count_0 == 0) && (_source_stream_matmul_23_source_21_pat_count_1 == 0)) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_cur_offset_2 <= _source_stream_matmul_23_source_21_pat_cur_offset_2 + _source_stream_matmul_23_source_21_pat_stride_buf_2;
        _source_stream_matmul_23_source_21_pat_count_2 <= _source_stream_matmul_23_source_21_pat_count_2 - 1;
      end 
      if((_stream_matmul_23_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_23_source_21_pat_count_0 == 0) && (_source_stream_matmul_23_source_21_pat_count_1 == 0)) && (_source_stream_matmul_23_source_21_pat_count_2 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_cur_offset_2 <= 0;
        _source_stream_matmul_23_source_21_pat_count_2 <= _source_stream_matmul_23_source_21_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_23_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_23_source_21_pat_count_0 == 0) && (_source_stream_matmul_23_source_21_pat_count_1 == 0) && (_source_stream_matmul_23_source_21_pat_count_2 == 0)) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_cur_offset_3 <= _source_stream_matmul_23_source_21_pat_cur_offset_3 + _source_stream_matmul_23_source_21_pat_stride_buf_3;
        _source_stream_matmul_23_source_21_pat_count_3 <= _source_stream_matmul_23_source_21_pat_count_3 - 1;
      end 
      if((_stream_matmul_23_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_23_source_21_pat_count_0 == 0) && (_source_stream_matmul_23_source_21_pat_count_1 == 0) && (_source_stream_matmul_23_source_21_pat_count_2 == 0)) && (_source_stream_matmul_23_source_21_pat_count_3 == 0) && _stream_matmul_23_stream_oready) begin
        _source_stream_matmul_23_source_21_pat_cur_offset_3 <= 0;
        _source_stream_matmul_23_source_21_pat_count_3 <= _source_stream_matmul_23_source_21_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_23_source_21_source_pat_fsm_3 == 1) && _stream_matmul_23_source_stop && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_21_source_ram_renable <= 0;
        _stream_matmul_23_source_21_idle <= 1;
      end 
      if((_stream_matmul_23_source_21_source_pat_fsm_3 == 2) && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_source_21_source_ram_renable <= 0;
        _stream_matmul_23_source_21_idle <= 1;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1412 <= _set_flag_1411;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1413 <= _tmp_1412;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1414 <= _tmp_1413;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1415 <= _tmp_1414;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1416 <= _tmp_1415;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1417 <= _tmp_1416;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1418 <= _tmp_1417;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1419 <= _tmp_1418;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1420 <= _tmp_1419;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1421 <= _tmp_1420;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1422 <= _tmp_1421;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1423 <= _tmp_1422;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1424 <= _tmp_1423;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1425 <= _tmp_1424;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1426 <= _tmp_1425;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1427 <= _tmp_1426;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1428 <= _tmp_1427;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1429 <= _tmp_1428;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1430 <= _tmp_1429;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1431 <= _tmp_1430;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1432 <= _tmp_1431;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1433 <= _tmp_1432;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1434 <= _tmp_1433;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1435 <= _tmp_1434;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1436 <= _tmp_1435;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1437 <= _tmp_1436;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1438 <= _tmp_1437;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1439 <= _tmp_1438;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1440 <= _tmp_1439;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1441 <= _tmp_1440;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1442 <= _tmp_1441;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1445 <= _tmp_1444;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1446 <= _tmp_1445;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1447 <= _tmp_1446;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1448 <= _tmp_1447;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1449 <= _tmp_1448;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1450 <= _tmp_1449;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1451 <= _tmp_1450;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1452 <= _tmp_1451;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1453 <= _tmp_1452;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1454 <= _tmp_1453;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1455 <= _tmp_1454;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1456 <= _tmp_1455;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1457 <= _tmp_1456;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1458 <= _tmp_1457;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1459 <= _tmp_1458;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1460 <= _tmp_1459;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1461 <= _tmp_1460;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1462 <= _tmp_1461;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1463 <= _tmp_1462;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1464 <= _tmp_1463;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1465 <= _tmp_1464;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1466 <= _tmp_1465;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1467 <= _tmp_1466;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1468 <= _tmp_1467;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1469 <= _tmp_1468;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1470 <= _tmp_1469;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1471 <= _tmp_1470;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1472 <= _tmp_1471;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1473 <= _tmp_1472;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1474 <= _tmp_1473;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1475 <= _tmp_1474;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1476 <= matmul_23_next_stream_num_ops;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1477 <= _tmp_1476;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1478 <= _tmp_1477;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1479 <= _tmp_1478;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1480 <= _tmp_1479;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1481 <= _tmp_1480;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1482 <= _tmp_1481;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1483 <= _tmp_1482;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1484 <= _tmp_1483;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1485 <= _tmp_1484;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1486 <= _tmp_1485;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1487 <= _tmp_1486;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1488 <= _tmp_1487;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1489 <= _tmp_1488;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1490 <= _tmp_1489;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1491 <= _tmp_1490;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1492 <= _tmp_1491;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1493 <= _tmp_1492;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1494 <= _tmp_1493;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1495 <= _tmp_1494;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1496 <= _tmp_1495;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1497 <= _tmp_1496;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1498 <= _tmp_1497;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1499 <= _tmp_1498;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1500 <= _tmp_1499;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1501 <= _tmp_1500;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1502 <= _tmp_1501;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1503 <= _tmp_1502;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1504 <= _tmp_1503;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1505 <= _tmp_1504;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1506 <= _tmp_1505;
      end 
      if(_tmp_1442) begin
        _stream_matmul_23_sink_26_sink_mode <= 5'b1;
        _stream_matmul_23_sink_26_sink_offset <= _tmp_1475;
        _stream_matmul_23_sink_26_sink_size <= _tmp_1506;
        _stream_matmul_23_sink_26_sink_stride <= 1;
      end 
      if(_tmp_1442) begin
        _stream_matmul_23_sink_26_sink_sel <= 5;
      end 
      if(_stream_matmul_23_sink_start && _stream_matmul_23_sink_26_sink_mode & 5'b1 && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_sink_26_sink_offset_buf <= _stream_matmul_23_sink_26_sink_offset;
        _stream_matmul_23_sink_26_sink_size_buf <= _stream_matmul_23_sink_26_sink_size;
        _stream_matmul_23_sink_26_sink_stride_buf <= _stream_matmul_23_sink_26_sink_stride;
      end 
      if((_stream_matmul_23_sink_26_sink_fsm_4 == 1) && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_sink_26_sink_waddr <= _stream_matmul_23_sink_26_sink_offset_buf - _stream_matmul_23_sink_26_sink_stride_buf;
        _stream_matmul_23_sink_26_sink_count <= _stream_matmul_23_sink_26_sink_size_buf;
      end 
      if((_stream_matmul_23_sink_26_sink_fsm_4 == 2) && stream_matmul_23_sink_27_data && _stream_matmul_23_stream_oready) begin
        _stream_matmul_23_sink_26_sink_waddr <= _stream_matmul_23_sink_26_sink_waddr + _stream_matmul_23_sink_26_sink_stride_buf;
        _stream_matmul_23_sink_26_sink_wdata <= stream_matmul_23_sink_26_data;
        _stream_matmul_23_sink_26_sink_wenable <= 1;
        _stream_matmul_23_sink_26_sink_count <= _stream_matmul_23_sink_26_sink_count - 1;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1519 <= _stream_matmul_23_source_start;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1520 <= _tmp_1519;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1521 <= _tmp_1520;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1522 <= _stream_matmul_23_source_start;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1523 <= _tmp_1522;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1524 <= _tmp_1523;
      end 
      if(_stream_matmul_23_stream_oready && _tmp_1524) begin
        __variable_wdata_961 <= 1;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1525 <= _stream_matmul_23_source_start;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1526 <= _tmp_1525;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1527 <= _tmp_1526;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1528 <= _tmp_1527;
      end 
      if(_stream_matmul_23_stream_oready && _tmp_1528) begin
        __variable_wdata_961 <= 0;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1531 <= _tmp_1530;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1534 <= _tmp_1533;
      end 
      if(_stream_matmul_23_stream_oready && _tmp_1534) begin
        __variable_wdata_961 <= 1;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1535 <= _stream_matmul_23_source_start;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1536 <= _tmp_1535;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1537 <= _tmp_1536;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1538 <= _tmp_1537;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1539 <= _tmp_1538;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1540 <= _tmp_1539;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1541 <= _tmp_1540;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1542 <= _tmp_1541;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1543 <= _tmp_1542;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1544 <= _tmp_1543;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1545 <= _tmp_1544;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1546 <= _tmp_1545;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1547 <= _tmp_1546;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1548 <= _tmp_1547;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1549 <= _tmp_1548;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1550 <= _tmp_1549;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1551 <= _tmp_1550;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1552 <= _tmp_1551;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1553 <= _tmp_1552;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1554 <= _tmp_1553;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1555 <= _tmp_1554;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1556 <= _tmp_1555;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1557 <= _tmp_1556;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1558 <= _tmp_1557;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1559 <= _tmp_1558;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1560 <= _tmp_1559;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1561 <= _tmp_1560;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1562 <= _tmp_1561;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1563 <= _tmp_1562;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1564 <= _tmp_1563;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1565 <= _tmp_1564;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1566 <= _stream_matmul_23_source_stop;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1567 <= _tmp_1566;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1568 <= _tmp_1567;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1569 <= _tmp_1568;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1570 <= _tmp_1569;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1571 <= _tmp_1570;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1572 <= _tmp_1571;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1573 <= _tmp_1572;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1574 <= _tmp_1573;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1575 <= _tmp_1574;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1576 <= _tmp_1575;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1577 <= _tmp_1576;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1578 <= _tmp_1577;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1579 <= _tmp_1578;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1580 <= _tmp_1579;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1581 <= _tmp_1580;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1582 <= _tmp_1581;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1583 <= _tmp_1582;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1584 <= _tmp_1583;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1585 <= _tmp_1584;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1586 <= _tmp_1585;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1587 <= _tmp_1586;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1588 <= _tmp_1587;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1589 <= _tmp_1588;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1590 <= _tmp_1589;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1591 <= _tmp_1590;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1592 <= _tmp_1591;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1593 <= _tmp_1592;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1594 <= _tmp_1593;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1595 <= _tmp_1594;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1596 <= _tmp_1595;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1597 <= _stream_matmul_23_source_busy;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1598 <= _tmp_1597;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1599 <= _tmp_1598;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1600 <= _tmp_1599;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1601 <= _tmp_1600;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1602 <= _tmp_1601;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1603 <= _tmp_1602;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1604 <= _tmp_1603;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1605 <= _tmp_1604;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1606 <= _tmp_1605;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1607 <= _tmp_1606;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1608 <= _tmp_1607;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1609 <= _tmp_1608;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1610 <= _tmp_1609;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1611 <= _tmp_1610;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1612 <= _tmp_1611;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1613 <= _tmp_1612;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1614 <= _tmp_1613;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1615 <= _tmp_1614;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1616 <= _tmp_1615;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1617 <= _tmp_1616;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1618 <= _tmp_1617;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1619 <= _tmp_1618;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1620 <= _tmp_1619;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1621 <= _tmp_1620;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1622 <= _tmp_1621;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1623 <= _tmp_1622;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1624 <= _tmp_1623;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1625 <= _tmp_1624;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1626 <= _tmp_1625;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1627 <= _tmp_1626;
      end 
      if(_stream_matmul_23_stream_oready) begin
        _tmp_1628 <= _stream_matmul_23_sink_busy;
      end 
      if(!_stream_matmul_23_sink_busy && _tmp_1628) begin
        _stream_matmul_23_busy_reg <= 0;
      end 
      if(_stream_matmul_23_source_busy) begin
        _stream_matmul_23_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_matmul_23_fsm_1 = 1;
  localparam _stream_matmul_23_fsm_2 = 2;
  localparam _stream_matmul_23_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_23_fsm <= _stream_matmul_23_fsm_init;
      _stream_matmul_23_source_start <= 0;
      _stream_matmul_23_source_busy <= 0;
      _stream_matmul_23_stream_ivalid <= 0;
    end else begin
      if(_stream_matmul_23_stream_oready && _tmp_1521) begin
        _stream_matmul_23_stream_ivalid <= 1;
      end 
      if(_stream_matmul_23_stream_oready && _tmp_1531) begin
        _stream_matmul_23_stream_ivalid <= 0;
      end 
      case(_stream_matmul_23_fsm)
        _stream_matmul_23_fsm_init: begin
          if(_stream_matmul_23_run_flag) begin
            _stream_matmul_23_source_start <= 1;
          end 
          if(_stream_matmul_23_run_flag) begin
            _stream_matmul_23_fsm <= _stream_matmul_23_fsm_1;
          end 
        end
        _stream_matmul_23_fsm_1: begin
          if(_stream_matmul_23_source_start && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_start <= 0;
            _stream_matmul_23_source_busy <= 1;
          end 
          if(_stream_matmul_23_source_start && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_fsm <= _stream_matmul_23_fsm_2;
          end 
        end
        _stream_matmul_23_fsm_2: begin
          if(_stream_matmul_23_stream_oready) begin
            _stream_matmul_23_fsm <= _stream_matmul_23_fsm_3;
          end 
        end
        _stream_matmul_23_fsm_3: begin
          if(_stream_matmul_23_stream_oready && (_stream_matmul_23_source_11_idle && _stream_matmul_23_source_13_idle && _stream_matmul_23_source_15_idle && _stream_matmul_23_source_20_idle && _stream_matmul_23_source_21_idle && _stream_matmul_23_source_7_idle && _stream_matmul_23_source_9_idle && (_stream_matmul_23_fsm == 3))) begin
            _stream_matmul_23_source_busy <= 0;
          end 
          if(_stream_matmul_23_stream_oready && (_stream_matmul_23_source_11_idle && _stream_matmul_23_source_13_idle && _stream_matmul_23_source_15_idle && _stream_matmul_23_source_20_idle && _stream_matmul_23_source_21_idle && _stream_matmul_23_source_7_idle && _stream_matmul_23_source_9_idle && (_stream_matmul_23_fsm == 3)) && _stream_matmul_23_run_flag) begin
            _stream_matmul_23_source_start <= 1;
          end 
          if(_stream_matmul_23_stream_oready && (_stream_matmul_23_source_11_idle && _stream_matmul_23_source_13_idle && _stream_matmul_23_source_15_idle && _stream_matmul_23_source_20_idle && _stream_matmul_23_source_21_idle && _stream_matmul_23_source_7_idle && _stream_matmul_23_source_9_idle && (_stream_matmul_23_fsm == 3))) begin
            _stream_matmul_23_fsm <= _stream_matmul_23_fsm_init;
          end 
          if(_stream_matmul_23_stream_oready && (_stream_matmul_23_source_11_idle && _stream_matmul_23_source_13_idle && _stream_matmul_23_source_15_idle && _stream_matmul_23_source_20_idle && _stream_matmul_23_source_21_idle && _stream_matmul_23_source_7_idle && _stream_matmul_23_source_9_idle && (_stream_matmul_23_fsm == 3)) && _stream_matmul_23_run_flag) begin
            _stream_matmul_23_fsm <= _stream_matmul_23_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_33_source_7_source_ram_renable <= 0;
      _stream_matmul_33_source_7_source_fifo_deq <= 0;
      _stream_matmul_33_source_7_idle <= 1;
      _stream_matmul_33_source_9_source_ram_renable <= 0;
      _stream_matmul_33_source_9_source_fifo_deq <= 0;
      _stream_matmul_33_source_9_idle <= 1;
      _stream_matmul_33_source_11_source_ram_renable <= 0;
      _stream_matmul_33_source_11_source_fifo_deq <= 0;
      _stream_matmul_33_source_11_idle <= 1;
      _stream_matmul_33_source_13_source_ram_renable <= 0;
      _stream_matmul_33_source_13_source_fifo_deq <= 0;
      _stream_matmul_33_source_13_idle <= 1;
      _stream_matmul_33_source_15_source_ram_renable <= 0;
      _stream_matmul_33_source_15_source_fifo_deq <= 0;
      _stream_matmul_33_source_15_idle <= 1;
      _stream_matmul_33_source_20_source_ram_renable <= 0;
      _stream_matmul_33_source_20_source_fifo_deq <= 0;
      _stream_matmul_33_source_20_idle <= 1;
      _stream_matmul_33_source_21_source_ram_renable <= 0;
      _stream_matmul_33_source_21_source_fifo_deq <= 0;
      _stream_matmul_33_source_21_idle <= 1;
      _stream_matmul_33_source_22_source_ram_renable <= 0;
      _stream_matmul_33_source_22_source_fifo_deq <= 0;
      _stream_matmul_33_source_22_idle <= 1;
      _stream_matmul_33_sink_33_sink_wenable <= 0;
      _stream_matmul_33_sink_33_sink_fifo_enq <= 0;
      _stream_matmul_33_sink_34_sink_wenable <= 0;
      _stream_matmul_33_sink_34_sink_fifo_enq <= 0;
      __stream_matmul_33_stream_ivalid_1 <= 0;
      __stream_matmul_33_stream_ivalid_2 <= 0;
      __stream_matmul_33_stream_ivalid_3 <= 0;
      __stream_matmul_33_stream_ivalid_4 <= 0;
      __stream_matmul_33_stream_ivalid_5 <= 0;
      __stream_matmul_33_stream_ivalid_6 <= 0;
      __stream_matmul_33_stream_ivalid_7 <= 0;
      __stream_matmul_33_stream_ivalid_8 <= 0;
      __stream_matmul_33_stream_ivalid_9 <= 0;
      __stream_matmul_33_stream_ivalid_10 <= 0;
      __stream_matmul_33_stream_ivalid_11 <= 0;
      __stream_matmul_33_stream_ivalid_12 <= 0;
      __stream_matmul_33_stream_ivalid_13 <= 0;
      __stream_matmul_33_stream_ivalid_14 <= 0;
      __stream_matmul_33_stream_ivalid_15 <= 0;
      __stream_matmul_33_stream_ivalid_16 <= 0;
      __stream_matmul_33_stream_ivalid_17 <= 0;
      __stream_matmul_33_stream_ivalid_18 <= 0;
      __stream_matmul_33_stream_ivalid_19 <= 0;
      __stream_matmul_33_stream_ivalid_20 <= 0;
      __stream_matmul_33_stream_ivalid_21 <= 0;
      __stream_matmul_33_stream_ivalid_22 <= 0;
      __stream_matmul_33_stream_ivalid_23 <= 0;
      __stream_matmul_33_stream_ivalid_24 <= 0;
      __stream_matmul_33_stream_ivalid_25 <= 0;
      __stream_matmul_33_stream_ivalid_26 <= 0;
      __stream_matmul_33_stream_ivalid_27 <= 0;
      __stream_matmul_33_stream_ivalid_28 <= 0;
      __stream_matmul_33_stream_ivalid_29 <= 0;
      __stream_matmul_33_stream_ivalid_30 <= 0;
      _counter_data_1058 <= 1'sd0;
      _counter_count_1058 <= 1'sd0;
      _minus_data_1063 <= 0;
      _minus_data_1069 <= 0;
      _eq_data_1138 <= 0;
      _eq_data_1142 <= 0;
      _plus_data_1189 <= 0;
      _plus_data_1194 <= 0;
      _plus_data_1199 <= 0;
      _plus_data_1204 <= 0;
      _plus_data_1210 <= 0;
      _plus_data_1215 <= 0;
      _plus_data_1231 <= 0;
      _plus_data_1250 <= 0;
      __delay_data_1501_pointer_1061 <= 0;
      __delay_data_1503__variable_1137 <= 0;
      __delay_data_1506_pointer_1184 <= 0;
      __delay_data_1509_reinterpretcast_1163 <= 0;
      __delay_data_1514_pointer_1067 <= 0;
      __delay_data_1518_reinterpretcast_1167 <= 0;
      __delay_data_1523__variable_1057 <= 0;
      __delay_data_1550__variable_1052 <= 0;
      __delay_data_1564_reinterpretcast_1175 <= 0;
      __delay_data_1569_reinterpretcast_1179 <= 0;
      __delay_data_1587_cond_1084 <= 0;
      __delay_data_1607_cond_1096 <= 0;
      __delay_data_1648_cond_1083 <= 0;
      __delay_data_1668_cond_1095 <= 0;
      _eq_data_1065 <= 0;
      _eq_data_1071 <= 0;
      __delay_data_1502__delay_1501_pointer_1061 <= 0;
      __delay_data_1504_reinterpretcast_1149 <= 0;
      __delay_data_1507__delay_1506_pointer_1184 <= 0;
      __delay_data_1510__delay_1509_reinterpretcast_1163 <= 0;
      __delay_data_1512_plus_1189 <= 0;
      __delay_data_1515__delay_1514_pointer_1067 <= 0;
      __delay_data_1516_reinterpretcast_1153 <= 0;
      __delay_data_1519__delay_1518_reinterpretcast_1167 <= 0;
      __delay_data_1521_plus_1194 <= 0;
      __delay_data_1524__delay_1523__variable_1057 <= 0;
      __delay_data_1537_plus_1199 <= 0;
      __delay_data_1551__delay_1550__variable_1052 <= 0;
      __delay_data_1565__delay_1564_reinterpretcast_1175 <= 0;
      __delay_data_1567_plus_1210 <= 0;
      __delay_data_1570__delay_1569_reinterpretcast_1179 <= 0;
      __delay_data_1572_plus_1215 <= 0;
      __delay_data_1574_plus_1231 <= 0;
      __delay_data_1588__delay_1587_cond_1084 <= 0;
      __delay_data_1608__delay_1607_cond_1096 <= 0;
      __delay_data_1628_plus_1250 <= 0;
      __delay_data_1649__delay_1648_cond_1083 <= 0;
      __delay_data_1669__delay_1668_cond_1095 <= 0;
      __delay_data_1689_plus_1204 <= 0;
      _land_data_1066 <= 0;
      _land_data_1072 <= 0;
      __delay_data_1505__delay_1504_reinterpretcast_1149 <= 0;
      __delay_data_1508__delay_1507__delay_1506_pointer_1184 <= 0;
      __delay_data_1511__delay_1510__delay_1509_reinterpretcast_1163 <= 0;
      __delay_data_1513__delay_1512_plus_1189 <= 0;
      __delay_data_1517__delay_1516_reinterpretcast_1153 <= 0;
      __delay_data_1520__delay_1519__delay_1518_reinterpretcast_1167 <= 0;
      __delay_data_1522__delay_1521_plus_1194 <= 0;
      __delay_data_1525__delay_1524__delay_1523__variable_1057 <= 0;
      __delay_data_1538__delay_1537_plus_1199 <= 0;
      __delay_data_1552__delay_1551__delay_1550__variable_1052 <= 0;
      __delay_data_1566__delay_1565__delay_1564_reinterpretcast_1175 <= 0;
      __delay_data_1568__delay_1567_plus_1210 <= 0;
      __delay_data_1571__delay_1570__delay_1569_reinterpretcast_1179 <= 0;
      __delay_data_1573__delay_1572_plus_1215 <= 0;
      __delay_data_1575__delay_1574_plus_1231 <= 0;
      __delay_data_1589__delay_1588__delay_1587_cond_1084 <= 0;
      __delay_data_1609__delay_1608__delay_1607_cond_1096 <= 0;
      __delay_data_1629__delay_1628_plus_1250 <= 0;
      __delay_data_1650__delay_1649__delay_1648_cond_1083 <= 0;
      __delay_data_1670__delay_1669__delay_1668_cond_1095 <= 0;
      __delay_data_1690__delay_1689_plus_1204 <= 0;
      __delay_data_1526__delay_1525__delay_1524____variable_1057 <= 0;
      __delay_data_1539__delay_1538__delay_1537_plus_1199 <= 0;
      __delay_data_1553__delay_1552__delay_1551____variable_1052 <= 0;
      __delay_data_1576__delay_1575__delay_1574_plus_1231 <= 0;
      __delay_data_1590__delay_1589__delay_1588___cond_1084 <= 0;
      __delay_data_1610__delay_1609__delay_1608___cond_1096 <= 0;
      __delay_data_1630__delay_1629__delay_1628_plus_1250 <= 0;
      __delay_data_1651__delay_1650__delay_1649___cond_1083 <= 0;
      __delay_data_1671__delay_1670__delay_1669___cond_1095 <= 0;
      __delay_data_1691__delay_1690__delay_1689_plus_1204 <= 0;
      __delay_data_1527__delay_1526__delay_1525____variable_1057 <= 0;
      __delay_data_1540__delay_1539__delay_1538___plus_1199 <= 0;
      __delay_data_1554__delay_1553__delay_1552____variable_1052 <= 0;
      __delay_data_1577__delay_1576__delay_1575___plus_1231 <= 0;
      __delay_data_1591__delay_1590__delay_1589___cond_1084 <= 0;
      __delay_data_1611__delay_1610__delay_1609___cond_1096 <= 0;
      __delay_data_1631__delay_1630__delay_1629___plus_1250 <= 0;
      __delay_data_1652__delay_1651__delay_1650___cond_1083 <= 0;
      __delay_data_1672__delay_1671__delay_1670___cond_1095 <= 0;
      __delay_data_1692__delay_1691__delay_1690___plus_1204 <= 0;
      __delay_data_1528__delay_1527__delay_1526____variable_1057 <= 0;
      __delay_data_1541__delay_1540__delay_1539___plus_1199 <= 0;
      __delay_data_1555__delay_1554__delay_1553____variable_1052 <= 0;
      __delay_data_1578__delay_1577__delay_1576___plus_1231 <= 0;
      __delay_data_1592__delay_1591__delay_1590___cond_1084 <= 0;
      __delay_data_1612__delay_1611__delay_1610___cond_1096 <= 0;
      __delay_data_1632__delay_1631__delay_1630___plus_1250 <= 0;
      __delay_data_1653__delay_1652__delay_1651___cond_1083 <= 0;
      __delay_data_1673__delay_1672__delay_1671___cond_1095 <= 0;
      __delay_data_1693__delay_1692__delay_1691___plus_1204 <= 0;
      __delay_data_1529__delay_1528__delay_1527____variable_1057 <= 0;
      __delay_data_1542__delay_1541__delay_1540___plus_1199 <= 0;
      __delay_data_1556__delay_1555__delay_1554____variable_1052 <= 0;
      __delay_data_1579__delay_1578__delay_1577___plus_1231 <= 0;
      __delay_data_1593__delay_1592__delay_1591___cond_1084 <= 0;
      __delay_data_1613__delay_1612__delay_1611___cond_1096 <= 0;
      __delay_data_1633__delay_1632__delay_1631___plus_1250 <= 0;
      __delay_data_1654__delay_1653__delay_1652___cond_1083 <= 0;
      __delay_data_1674__delay_1673__delay_1672___cond_1095 <= 0;
      __delay_data_1694__delay_1693__delay_1692___plus_1204 <= 0;
      __delay_data_1530__delay_1529__delay_1528____variable_1057 <= 0;
      __delay_data_1543__delay_1542__delay_1541___plus_1199 <= 0;
      __delay_data_1557__delay_1556__delay_1555____variable_1052 <= 0;
      __delay_data_1580__delay_1579__delay_1578___plus_1231 <= 0;
      __delay_data_1594__delay_1593__delay_1592___cond_1084 <= 0;
      __delay_data_1614__delay_1613__delay_1612___cond_1096 <= 0;
      __delay_data_1634__delay_1633__delay_1632___plus_1250 <= 0;
      __delay_data_1655__delay_1654__delay_1653___cond_1083 <= 0;
      __delay_data_1675__delay_1674__delay_1673___cond_1095 <= 0;
      __delay_data_1695__delay_1694__delay_1693___plus_1204 <= 0;
      __delay_data_1531__delay_1530__delay_1529____variable_1057 <= 0;
      __delay_data_1544__delay_1543__delay_1542___plus_1199 <= 0;
      __delay_data_1558__delay_1557__delay_1556____variable_1052 <= 0;
      __delay_data_1581__delay_1580__delay_1579___plus_1231 <= 0;
      __delay_data_1595__delay_1594__delay_1593___cond_1084 <= 0;
      __delay_data_1615__delay_1614__delay_1613___cond_1096 <= 0;
      __delay_data_1635__delay_1634__delay_1633___plus_1250 <= 0;
      __delay_data_1656__delay_1655__delay_1654___cond_1083 <= 0;
      __delay_data_1676__delay_1675__delay_1674___cond_1095 <= 0;
      __delay_data_1696__delay_1695__delay_1694___plus_1204 <= 0;
      __delay_data_1532__delay_1531__delay_1530____variable_1057 <= 0;
      __delay_data_1545__delay_1544__delay_1543___plus_1199 <= 0;
      __delay_data_1559__delay_1558__delay_1557____variable_1052 <= 0;
      __delay_data_1582__delay_1581__delay_1580___plus_1231 <= 0;
      __delay_data_1596__delay_1595__delay_1594___cond_1084 <= 0;
      __delay_data_1616__delay_1615__delay_1614___cond_1096 <= 0;
      __delay_data_1636__delay_1635__delay_1634___plus_1250 <= 0;
      __delay_data_1657__delay_1656__delay_1655___cond_1083 <= 0;
      __delay_data_1677__delay_1676__delay_1675___cond_1095 <= 0;
      __delay_data_1697__delay_1696__delay_1695___plus_1204 <= 0;
      __delay_data_1533__delay_1532__delay_1531____variable_1057 <= 0;
      __delay_data_1546__delay_1545__delay_1544___plus_1199 <= 0;
      __delay_data_1560__delay_1559__delay_1558____variable_1052 <= 0;
      __delay_data_1583__delay_1582__delay_1581___plus_1231 <= 0;
      __delay_data_1597__delay_1596__delay_1595___cond_1084 <= 0;
      __delay_data_1617__delay_1616__delay_1615___cond_1096 <= 0;
      __delay_data_1637__delay_1636__delay_1635___plus_1250 <= 0;
      __delay_data_1658__delay_1657__delay_1656___cond_1083 <= 0;
      __delay_data_1678__delay_1677__delay_1676___cond_1095 <= 0;
      __delay_data_1698__delay_1697__delay_1696___plus_1204 <= 0;
      __delay_data_1534__delay_1533__delay_1532____variable_1057 <= 0;
      __delay_data_1547__delay_1546__delay_1545___plus_1199 <= 0;
      __delay_data_1561__delay_1560__delay_1559____variable_1052 <= 0;
      __delay_data_1584__delay_1583__delay_1582___plus_1231 <= 0;
      __delay_data_1598__delay_1597__delay_1596___cond_1084 <= 0;
      __delay_data_1618__delay_1617__delay_1616___cond_1096 <= 0;
      __delay_data_1638__delay_1637__delay_1636___plus_1250 <= 0;
      __delay_data_1659__delay_1658__delay_1657___cond_1083 <= 0;
      __delay_data_1679__delay_1678__delay_1677___cond_1095 <= 0;
      __delay_data_1699__delay_1698__delay_1697___plus_1204 <= 0;
      __delay_data_1535__delay_1534__delay_1533____variable_1057 <= 0;
      __delay_data_1548__delay_1547__delay_1546___plus_1199 <= 0;
      __delay_data_1562__delay_1561__delay_1560____variable_1052 <= 0;
      __delay_data_1585__delay_1584__delay_1583___plus_1231 <= 0;
      __delay_data_1599__delay_1598__delay_1597___cond_1084 <= 0;
      __delay_data_1619__delay_1618__delay_1617___cond_1096 <= 0;
      __delay_data_1639__delay_1638__delay_1637___plus_1250 <= 0;
      __delay_data_1660__delay_1659__delay_1658___cond_1083 <= 0;
      __delay_data_1680__delay_1679__delay_1678___cond_1095 <= 0;
      __delay_data_1700__delay_1699__delay_1698___plus_1204 <= 0;
      __delay_data_1536__delay_1535__delay_1534____variable_1057 <= 0;
      __delay_data_1549__delay_1548__delay_1547___plus_1199 <= 0;
      __delay_data_1563__delay_1562__delay_1561____variable_1052 <= 0;
      __delay_data_1586__delay_1585__delay_1584___plus_1231 <= 0;
      __delay_data_1600__delay_1599__delay_1598___cond_1084 <= 0;
      __delay_data_1620__delay_1619__delay_1618___cond_1096 <= 0;
      __delay_data_1640__delay_1639__delay_1638___plus_1250 <= 0;
      __delay_data_1661__delay_1660__delay_1659___cond_1083 <= 0;
      __delay_data_1681__delay_1680__delay_1679___cond_1095 <= 0;
      __delay_data_1701__delay_1700__delay_1699___plus_1204 <= 0;
      __delay_data_1601__delay_1600__delay_1599___cond_1084 <= 0;
      __delay_data_1621__delay_1620__delay_1619___cond_1096 <= 0;
      __delay_data_1641__delay_1640__delay_1639___plus_1250 <= 0;
      __delay_data_1662__delay_1661__delay_1660___cond_1083 <= 0;
      __delay_data_1682__delay_1681__delay_1680___cond_1095 <= 0;
      __delay_data_1702__delay_1701__delay_1700___plus_1204 <= 0;
      __delay_data_1602__delay_1601__delay_1600___cond_1084 <= 0;
      __delay_data_1622__delay_1621__delay_1620___cond_1096 <= 0;
      __delay_data_1642__delay_1641__delay_1640___plus_1250 <= 0;
      __delay_data_1663__delay_1662__delay_1661___cond_1083 <= 0;
      __delay_data_1683__delay_1682__delay_1681___cond_1095 <= 0;
      __delay_data_1703__delay_1702__delay_1701___plus_1204 <= 0;
      __delay_data_1603__delay_1602__delay_1601___cond_1084 <= 0;
      __delay_data_1623__delay_1622__delay_1621___cond_1096 <= 0;
      __delay_data_1643__delay_1642__delay_1641___plus_1250 <= 0;
      __delay_data_1664__delay_1663__delay_1662___cond_1083 <= 0;
      __delay_data_1684__delay_1683__delay_1682___cond_1095 <= 0;
      __delay_data_1704__delay_1703__delay_1702___plus_1204 <= 0;
      __delay_data_1604__delay_1603__delay_1602___cond_1084 <= 0;
      __delay_data_1624__delay_1623__delay_1622___cond_1096 <= 0;
      __delay_data_1644__delay_1643__delay_1642___plus_1250 <= 0;
      __delay_data_1665__delay_1664__delay_1663___cond_1083 <= 0;
      __delay_data_1685__delay_1684__delay_1683___cond_1095 <= 0;
      __delay_data_1705__delay_1704__delay_1703___plus_1204 <= 0;
      __delay_data_1605__delay_1604__delay_1603___cond_1084 <= 0;
      __delay_data_1625__delay_1624__delay_1623___cond_1096 <= 0;
      __delay_data_1645__delay_1644__delay_1643___plus_1250 <= 0;
      __delay_data_1666__delay_1665__delay_1664___cond_1083 <= 0;
      __delay_data_1686__delay_1685__delay_1684___cond_1095 <= 0;
      __delay_data_1706__delay_1705__delay_1704___plus_1204 <= 0;
      __delay_data_1606__delay_1605__delay_1604___cond_1084 <= 0;
      __delay_data_1626__delay_1625__delay_1624___cond_1096 <= 0;
      __delay_data_1646__delay_1645__delay_1644___plus_1250 <= 0;
      __delay_data_1667__delay_1666__delay_1665___cond_1083 <= 0;
      __delay_data_1687__delay_1686__delay_1685___cond_1095 <= 0;
      __delay_data_1707__delay_1706__delay_1705___plus_1204 <= 0;
      _plus_data_1202 <= 0;
      _plus_data_1234 <= 0;
      __delay_data_1627__delay_1626__delay_1625___cond_1096 <= 0;
      __delay_data_1647__delay_1646__delay_1645___plus_1250 <= 0;
      __delay_data_1688__delay_1687__delay_1686___cond_1095 <= 0;
      __delay_data_1708__delay_1707__delay_1706___plus_1204 <= 0;
      __delay_data_1709__substreamoutput_1201 <= 0;
      __delay_data_1710__delay_1709__substreamoutput_1201 <= 0;
      __delay_data_1711__delay_1710____substreamoutput_1201 <= 0;
      __delay_data_1712__delay_1711____substreamoutput_1201 <= 0;
      __delay_data_1713__delay_1712____substreamoutput_1201 <= 0;
      __delay_data_1714__delay_1713____substreamoutput_1201 <= 0;
      __delay_data_1715__delay_1714____substreamoutput_1201 <= 0;
      __delay_data_1716__delay_1715____substreamoutput_1201 <= 0;
      __delay_data_1717__delay_1716____substreamoutput_1201 <= 0;
      __delay_data_1718__delay_1717____substreamoutput_1201 <= 0;
      _stream_matmul_33_parameter_0_next_parameter_data <= 0;
      __variable_wdata_1052 <= 0;
      _stream_matmul_33_parameter_1_next_parameter_data <= 0;
      __variable_wdata_1053 <= 0;
      _stream_matmul_33_parameter_2_next_parameter_data <= 0;
      __variable_wdata_1054 <= 0;
      _stream_matmul_33_parameter_3_next_parameter_data <= 0;
      __variable_wdata_1055 <= 0;
      _stream_matmul_33_parameter_4_next_parameter_data <= 0;
      __variable_wdata_1056 <= 0;
      _stream_matmul_33_parameter_6_next_parameter_data <= 0;
      __variable_wdata_1073 <= 0;
      _stream_matmul_33_source_7_source_mode <= 5'b0;
      _stream_matmul_33_source_7_source_offset <= 0;
      _source_stream_matmul_33_source_7_pat_size_0 <= 0;
      _source_stream_matmul_33_source_7_pat_stride_0 <= 0;
      _source_stream_matmul_33_source_7_pat_size_1 <= 0;
      _source_stream_matmul_33_source_7_pat_stride_1 <= 0;
      _source_stream_matmul_33_source_7_pat_size_2 <= 0;
      _source_stream_matmul_33_source_7_pat_stride_2 <= 0;
      _source_stream_matmul_33_source_7_pat_size_3 <= 0;
      _source_stream_matmul_33_source_7_pat_stride_3 <= 0;
      _stream_matmul_33_source_7_source_sel <= 0;
      _stream_matmul_33_source_7_source_offset_buf <= 0;
      _source_stream_matmul_33_source_7_pat_cur_offset_0 <= 0;
      _source_stream_matmul_33_source_7_pat_cur_offset_1 <= 0;
      _source_stream_matmul_33_source_7_pat_cur_offset_2 <= 0;
      _source_stream_matmul_33_source_7_pat_cur_offset_3 <= 0;
      _source_stream_matmul_33_source_7_pat_count_0 <= 0;
      _source_stream_matmul_33_source_7_pat_count_1 <= 0;
      _source_stream_matmul_33_source_7_pat_count_2 <= 0;
      _source_stream_matmul_33_source_7_pat_count_3 <= 0;
      _source_stream_matmul_33_source_7_pat_size_buf_0 <= 0;
      _source_stream_matmul_33_source_7_pat_size_buf_1 <= 0;
      _source_stream_matmul_33_source_7_pat_size_buf_2 <= 0;
      _source_stream_matmul_33_source_7_pat_size_buf_3 <= 0;
      _source_stream_matmul_33_source_7_pat_stride_buf_0 <= 0;
      _source_stream_matmul_33_source_7_pat_stride_buf_1 <= 0;
      _source_stream_matmul_33_source_7_pat_stride_buf_2 <= 0;
      _source_stream_matmul_33_source_7_pat_stride_buf_3 <= 0;
      __variable_wdata_1074 <= 0;
      _stream_matmul_33_source_7_source_ram_raddr <= 0;
      _stream_matmul_33_parameter_8_next_parameter_data <= 0;
      __variable_wdata_1085 <= 0;
      _stream_matmul_33_source_9_source_mode <= 5'b0;
      _stream_matmul_33_source_9_source_offset <= 0;
      _source_stream_matmul_33_source_9_pat_size_0 <= 0;
      _source_stream_matmul_33_source_9_pat_stride_0 <= 0;
      _source_stream_matmul_33_source_9_pat_size_1 <= 0;
      _source_stream_matmul_33_source_9_pat_stride_1 <= 0;
      _source_stream_matmul_33_source_9_pat_size_2 <= 0;
      _source_stream_matmul_33_source_9_pat_stride_2 <= 0;
      _source_stream_matmul_33_source_9_pat_size_3 <= 0;
      _source_stream_matmul_33_source_9_pat_stride_3 <= 0;
      _stream_matmul_33_source_9_source_sel <= 0;
      _stream_matmul_33_source_9_source_offset_buf <= 0;
      _source_stream_matmul_33_source_9_pat_cur_offset_0 <= 0;
      _source_stream_matmul_33_source_9_pat_cur_offset_1 <= 0;
      _source_stream_matmul_33_source_9_pat_cur_offset_2 <= 0;
      _source_stream_matmul_33_source_9_pat_cur_offset_3 <= 0;
      _source_stream_matmul_33_source_9_pat_count_0 <= 0;
      _source_stream_matmul_33_source_9_pat_count_1 <= 0;
      _source_stream_matmul_33_source_9_pat_count_2 <= 0;
      _source_stream_matmul_33_source_9_pat_count_3 <= 0;
      _source_stream_matmul_33_source_9_pat_size_buf_0 <= 0;
      _source_stream_matmul_33_source_9_pat_size_buf_1 <= 0;
      _source_stream_matmul_33_source_9_pat_size_buf_2 <= 0;
      _source_stream_matmul_33_source_9_pat_size_buf_3 <= 0;
      _source_stream_matmul_33_source_9_pat_stride_buf_0 <= 0;
      _source_stream_matmul_33_source_9_pat_stride_buf_1 <= 0;
      _source_stream_matmul_33_source_9_pat_stride_buf_2 <= 0;
      _source_stream_matmul_33_source_9_pat_stride_buf_3 <= 0;
      __variable_wdata_1086 <= 0;
      _stream_matmul_33_source_9_source_ram_raddr <= 0;
      _stream_matmul_33_parameter_10_next_parameter_data <= 0;
      __variable_wdata_1097 <= 0;
      _stream_matmul_33_source_11_source_mode <= 5'b0;
      _stream_matmul_33_source_11_source_empty_data <= 0;
      __variable_wdata_1098 <= 0;
      _stream_matmul_33_parameter_12_next_parameter_data <= 0;
      __variable_wdata_1109 <= 0;
      _stream_matmul_33_source_13_source_mode <= 5'b0;
      _stream_matmul_33_source_13_source_empty_data <= 0;
      __variable_wdata_1110 <= 0;
      _stream_matmul_33_parameter_14_next_parameter_data <= 0;
      __variable_wdata_1121 <= 0;
      _stream_matmul_33_source_15_source_mode <= 5'b0;
      _stream_matmul_33_source_15_source_empty_data <= 0;
      __variable_wdata_1122 <= 0;
      _stream_matmul_33_parameter_16_next_parameter_data <= 0;
      __variable_wdata_1133 <= 0;
      _stream_matmul_33_parameter_17_next_parameter_data <= 0;
      __variable_wdata_1134 <= 0;
      _stream_matmul_33_parameter_18_next_parameter_data <= 0;
      __variable_wdata_1135 <= 0;
      _stream_matmul_33_parameter_19_next_parameter_data <= 0;
      __variable_wdata_1136 <= 0;
      _stream_matmul_33_source_20_source_mode <= 5'b0;
      _stream_matmul_33_source_20_source_offset <= 0;
      _source_stream_matmul_33_source_20_pat_size_0 <= 0;
      _source_stream_matmul_33_source_20_pat_stride_0 <= 0;
      _source_stream_matmul_33_source_20_pat_size_1 <= 0;
      _source_stream_matmul_33_source_20_pat_stride_1 <= 0;
      _source_stream_matmul_33_source_20_pat_size_2 <= 0;
      _source_stream_matmul_33_source_20_pat_stride_2 <= 0;
      _source_stream_matmul_33_source_20_pat_size_3 <= 0;
      _source_stream_matmul_33_source_20_pat_stride_3 <= 0;
      _stream_matmul_33_source_20_source_sel <= 0;
      _stream_matmul_33_source_20_source_offset_buf <= 0;
      _source_stream_matmul_33_source_20_pat_cur_offset_0 <= 0;
      _source_stream_matmul_33_source_20_pat_cur_offset_1 <= 0;
      _source_stream_matmul_33_source_20_pat_cur_offset_2 <= 0;
      _source_stream_matmul_33_source_20_pat_cur_offset_3 <= 0;
      _source_stream_matmul_33_source_20_pat_count_0 <= 0;
      _source_stream_matmul_33_source_20_pat_count_1 <= 0;
      _source_stream_matmul_33_source_20_pat_count_2 <= 0;
      _source_stream_matmul_33_source_20_pat_count_3 <= 0;
      _source_stream_matmul_33_source_20_pat_size_buf_0 <= 0;
      _source_stream_matmul_33_source_20_pat_size_buf_1 <= 0;
      _source_stream_matmul_33_source_20_pat_size_buf_2 <= 0;
      _source_stream_matmul_33_source_20_pat_size_buf_3 <= 0;
      _source_stream_matmul_33_source_20_pat_stride_buf_0 <= 0;
      _source_stream_matmul_33_source_20_pat_stride_buf_1 <= 0;
      _source_stream_matmul_33_source_20_pat_stride_buf_2 <= 0;
      _source_stream_matmul_33_source_20_pat_stride_buf_3 <= 0;
      __variable_wdata_1137 <= 0;
      _stream_matmul_33_source_20_source_ram_raddr <= 0;
      _stream_matmul_33_source_21_source_mode <= 5'b0;
      _stream_matmul_33_source_21_source_offset <= 0;
      _source_stream_matmul_33_source_21_pat_size_0 <= 0;
      _source_stream_matmul_33_source_21_pat_stride_0 <= 0;
      _source_stream_matmul_33_source_21_pat_size_1 <= 0;
      _source_stream_matmul_33_source_21_pat_stride_1 <= 0;
      _source_stream_matmul_33_source_21_pat_size_2 <= 0;
      _source_stream_matmul_33_source_21_pat_stride_2 <= 0;
      _source_stream_matmul_33_source_21_pat_size_3 <= 0;
      _source_stream_matmul_33_source_21_pat_stride_3 <= 0;
      _stream_matmul_33_source_21_source_sel <= 0;
      _stream_matmul_33_source_21_source_offset_buf <= 0;
      _source_stream_matmul_33_source_21_pat_cur_offset_0 <= 0;
      _source_stream_matmul_33_source_21_pat_cur_offset_1 <= 0;
      _source_stream_matmul_33_source_21_pat_cur_offset_2 <= 0;
      _source_stream_matmul_33_source_21_pat_cur_offset_3 <= 0;
      _source_stream_matmul_33_source_21_pat_count_0 <= 0;
      _source_stream_matmul_33_source_21_pat_count_1 <= 0;
      _source_stream_matmul_33_source_21_pat_count_2 <= 0;
      _source_stream_matmul_33_source_21_pat_count_3 <= 0;
      _source_stream_matmul_33_source_21_pat_size_buf_0 <= 0;
      _source_stream_matmul_33_source_21_pat_size_buf_1 <= 0;
      _source_stream_matmul_33_source_21_pat_size_buf_2 <= 0;
      _source_stream_matmul_33_source_21_pat_size_buf_3 <= 0;
      _source_stream_matmul_33_source_21_pat_stride_buf_0 <= 0;
      _source_stream_matmul_33_source_21_pat_stride_buf_1 <= 0;
      _source_stream_matmul_33_source_21_pat_stride_buf_2 <= 0;
      _source_stream_matmul_33_source_21_pat_stride_buf_3 <= 0;
      __variable_wdata_1158 <= 0;
      _stream_matmul_33_source_21_source_ram_raddr <= 0;
      _stream_matmul_33_source_22_source_mode <= 5'b0;
      _stream_matmul_33_source_22_source_offset <= 0;
      _source_stream_matmul_33_source_22_pat_size_0 <= 0;
      _source_stream_matmul_33_source_22_pat_stride_0 <= 0;
      _source_stream_matmul_33_source_22_pat_size_1 <= 0;
      _source_stream_matmul_33_source_22_pat_stride_1 <= 0;
      _source_stream_matmul_33_source_22_pat_size_2 <= 0;
      _source_stream_matmul_33_source_22_pat_stride_2 <= 0;
      _source_stream_matmul_33_source_22_pat_size_3 <= 0;
      _source_stream_matmul_33_source_22_pat_stride_3 <= 0;
      _stream_matmul_33_source_22_source_sel <= 0;
      _stream_matmul_33_source_22_source_offset_buf <= 0;
      _source_stream_matmul_33_source_22_pat_cur_offset_0 <= 0;
      _source_stream_matmul_33_source_22_pat_cur_offset_1 <= 0;
      _source_stream_matmul_33_source_22_pat_cur_offset_2 <= 0;
      _source_stream_matmul_33_source_22_pat_cur_offset_3 <= 0;
      _source_stream_matmul_33_source_22_pat_count_0 <= 0;
      _source_stream_matmul_33_source_22_pat_count_1 <= 0;
      _source_stream_matmul_33_source_22_pat_count_2 <= 0;
      _source_stream_matmul_33_source_22_pat_count_3 <= 0;
      _source_stream_matmul_33_source_22_pat_size_buf_0 <= 0;
      _source_stream_matmul_33_source_22_pat_size_buf_1 <= 0;
      _source_stream_matmul_33_source_22_pat_size_buf_2 <= 0;
      _source_stream_matmul_33_source_22_pat_size_buf_3 <= 0;
      _source_stream_matmul_33_source_22_pat_stride_buf_0 <= 0;
      _source_stream_matmul_33_source_22_pat_stride_buf_1 <= 0;
      _source_stream_matmul_33_source_22_pat_stride_buf_2 <= 0;
      _source_stream_matmul_33_source_22_pat_stride_buf_3 <= 0;
      __variable_wdata_1159 <= 0;
      _stream_matmul_33_source_22_source_ram_raddr <= 0;
      _tmp_1703 <= 0;
      _tmp_1704 <= 0;
      _tmp_1705 <= 0;
      _tmp_1706 <= 0;
      _tmp_1707 <= 0;
      _tmp_1708 <= 0;
      _tmp_1709 <= 0;
      _tmp_1710 <= 0;
      _tmp_1711 <= 0;
      _tmp_1712 <= 0;
      _tmp_1713 <= 0;
      _tmp_1714 <= 0;
      _tmp_1715 <= 0;
      _tmp_1716 <= 0;
      _tmp_1717 <= 0;
      _tmp_1718 <= 0;
      _tmp_1719 <= 0;
      _tmp_1720 <= 0;
      _tmp_1721 <= 0;
      _tmp_1722 <= 0;
      _tmp_1723 <= 0;
      _tmp_1724 <= 0;
      _tmp_1725 <= 0;
      _tmp_1726 <= 0;
      _tmp_1727 <= 0;
      _tmp_1728 <= 0;
      _tmp_1729 <= 0;
      _tmp_1730 <= 0;
      _tmp_1731 <= 0;
      _tmp_1732 <= 0;
      _tmp_1733 <= 0;
      _tmp_1734 <= 0;
      _tmp_1737 <= 0;
      _tmp_1738 <= 0;
      _tmp_1739 <= 0;
      _tmp_1740 <= 0;
      _tmp_1741 <= 0;
      _tmp_1742 <= 0;
      _tmp_1743 <= 0;
      _tmp_1744 <= 0;
      _tmp_1745 <= 0;
      _tmp_1746 <= 0;
      _tmp_1747 <= 0;
      _tmp_1748 <= 0;
      _tmp_1749 <= 0;
      _tmp_1750 <= 0;
      _tmp_1751 <= 0;
      _tmp_1752 <= 0;
      _tmp_1753 <= 0;
      _tmp_1754 <= 0;
      _tmp_1755 <= 0;
      _tmp_1756 <= 0;
      _tmp_1757 <= 0;
      _tmp_1758 <= 0;
      _tmp_1759 <= 0;
      _tmp_1760 <= 0;
      _tmp_1761 <= 0;
      _tmp_1762 <= 0;
      _tmp_1763 <= 0;
      _tmp_1764 <= 0;
      _tmp_1765 <= 0;
      _tmp_1766 <= 0;
      _tmp_1767 <= 0;
      _tmp_1768 <= 0;
      _tmp_1769 <= 0;
      _tmp_1770 <= 0;
      _tmp_1771 <= 0;
      _tmp_1772 <= 0;
      _tmp_1773 <= 0;
      _tmp_1774 <= 0;
      _tmp_1775 <= 0;
      _tmp_1776 <= 0;
      _tmp_1777 <= 0;
      _tmp_1778 <= 0;
      _tmp_1779 <= 0;
      _tmp_1780 <= 0;
      _tmp_1781 <= 0;
      _tmp_1782 <= 0;
      _tmp_1783 <= 0;
      _tmp_1784 <= 0;
      _tmp_1785 <= 0;
      _tmp_1786 <= 0;
      _tmp_1787 <= 0;
      _tmp_1788 <= 0;
      _tmp_1789 <= 0;
      _tmp_1790 <= 0;
      _tmp_1791 <= 0;
      _tmp_1792 <= 0;
      _tmp_1793 <= 0;
      _tmp_1794 <= 0;
      _tmp_1795 <= 0;
      _tmp_1796 <= 0;
      _tmp_1797 <= 0;
      _tmp_1798 <= 0;
      _tmp_1799 <= 0;
      _tmp_1800 <= 0;
      _stream_matmul_33_sink_33_sink_mode <= 5'b0;
      _stream_matmul_33_sink_33_sink_offset <= 0;
      _stream_matmul_33_sink_33_sink_size <= 0;
      _stream_matmul_33_sink_33_sink_stride <= 0;
      _stream_matmul_33_sink_33_sink_sel <= 0;
      _stream_matmul_33_sink_33_sink_offset_buf <= 0;
      _stream_matmul_33_sink_33_sink_size_buf <= 0;
      _stream_matmul_33_sink_33_sink_stride_buf <= 0;
      _stream_matmul_33_sink_33_sink_waddr <= 0;
      _stream_matmul_33_sink_33_sink_count <= 0;
      _stream_matmul_33_sink_33_sink_wdata <= 0;
      _tmp_1894 <= 0;
      _tmp_1895 <= 0;
      _tmp_1896 <= 0;
      _tmp_1897 <= 0;
      _tmp_1898 <= 0;
      _tmp_1899 <= 0;
      __variable_wdata_1057 <= 0;
      _tmp_1900 <= 0;
      _tmp_1901 <= 0;
      _tmp_1902 <= 0;
      _tmp_1903 <= 0;
      _tmp_1906 <= 0;
      _tmp_1909 <= 0;
      _tmp_1910 <= 0;
      _tmp_1911 <= 0;
      _tmp_1912 <= 0;
      _tmp_1913 <= 0;
      _tmp_1914 <= 0;
      _tmp_1915 <= 0;
      _tmp_1916 <= 0;
      _tmp_1917 <= 0;
      _tmp_1918 <= 0;
      _tmp_1919 <= 0;
      _tmp_1920 <= 0;
      _tmp_1921 <= 0;
      _tmp_1922 <= 0;
      _tmp_1923 <= 0;
      _tmp_1924 <= 0;
      _tmp_1925 <= 0;
      _tmp_1926 <= 0;
      _tmp_1927 <= 0;
      _tmp_1928 <= 0;
      _tmp_1929 <= 0;
      _tmp_1930 <= 0;
      _tmp_1931 <= 0;
      _tmp_1932 <= 0;
      _tmp_1933 <= 0;
      _tmp_1934 <= 0;
      _tmp_1935 <= 0;
      _tmp_1936 <= 0;
      _tmp_1937 <= 0;
      _tmp_1938 <= 0;
      _tmp_1939 <= 0;
      _tmp_1940 <= 0;
      _tmp_1941 <= 0;
      _tmp_1942 <= 0;
      _tmp_1943 <= 0;
      _tmp_1944 <= 0;
      _tmp_1945 <= 0;
      _tmp_1946 <= 0;
      _tmp_1947 <= 0;
      _tmp_1948 <= 0;
      _tmp_1949 <= 0;
      _tmp_1950 <= 0;
      _tmp_1951 <= 0;
      _tmp_1952 <= 0;
      _tmp_1953 <= 0;
      _tmp_1954 <= 0;
      _tmp_1955 <= 0;
      _tmp_1956 <= 0;
      _tmp_1957 <= 0;
      _tmp_1958 <= 0;
      _tmp_1959 <= 0;
      _tmp_1960 <= 0;
      _tmp_1961 <= 0;
      _tmp_1962 <= 0;
      _tmp_1963 <= 0;
      _tmp_1964 <= 0;
      _tmp_1965 <= 0;
      _tmp_1966 <= 0;
      _tmp_1967 <= 0;
      _tmp_1968 <= 0;
      _tmp_1969 <= 0;
      _tmp_1970 <= 0;
      _tmp_1971 <= 0;
      _tmp_1972 <= 0;
      _tmp_1973 <= 0;
      _tmp_1974 <= 0;
      _tmp_1975 <= 0;
      _tmp_1976 <= 0;
      _tmp_1977 <= 0;
      _tmp_1978 <= 0;
      _tmp_1979 <= 0;
      _tmp_1980 <= 0;
      _tmp_1981 <= 0;
      _tmp_1982 <= 0;
      _tmp_1983 <= 0;
      _tmp_1984 <= 0;
      _tmp_1985 <= 0;
      _tmp_1986 <= 0;
      _tmp_1987 <= 0;
      _tmp_1988 <= 0;
      _tmp_1989 <= 0;
      _tmp_1990 <= 0;
      _tmp_1991 <= 0;
      _tmp_1992 <= 0;
      _tmp_1993 <= 0;
      _tmp_1994 <= 0;
      _tmp_1995 <= 0;
      _tmp_1996 <= 0;
      _tmp_1997 <= 0;
      _tmp_1998 <= 0;
      _tmp_1999 <= 0;
      _tmp_2000 <= 0;
      _tmp_2001 <= 0;
      _tmp_2002 <= 0;
      _tmp_2003 <= 0;
      _tmp_2004 <= 0;
      _tmp_2005 <= 0;
      _tmp_2006 <= 0;
      _stream_matmul_33_busy_reg <= 0;
    end else begin
      if(_stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_7_source_ram_renable <= 0;
        _stream_matmul_33_source_7_source_fifo_deq <= 0;
      end 
      _stream_matmul_33_source_7_idle <= _stream_matmul_33_source_7_idle;
      if(_stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_9_source_ram_renable <= 0;
        _stream_matmul_33_source_9_source_fifo_deq <= 0;
      end 
      _stream_matmul_33_source_9_idle <= _stream_matmul_33_source_9_idle;
      if(_stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_11_source_ram_renable <= 0;
        _stream_matmul_33_source_11_source_fifo_deq <= 0;
      end 
      _stream_matmul_33_source_11_idle <= _stream_matmul_33_source_11_idle;
      if(_stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_13_source_ram_renable <= 0;
        _stream_matmul_33_source_13_source_fifo_deq <= 0;
      end 
      _stream_matmul_33_source_13_idle <= _stream_matmul_33_source_13_idle;
      if(_stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_15_source_ram_renable <= 0;
        _stream_matmul_33_source_15_source_fifo_deq <= 0;
      end 
      _stream_matmul_33_source_15_idle <= _stream_matmul_33_source_15_idle;
      if(_stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_20_source_ram_renable <= 0;
        _stream_matmul_33_source_20_source_fifo_deq <= 0;
      end 
      _stream_matmul_33_source_20_idle <= _stream_matmul_33_source_20_idle;
      if(_stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_21_source_ram_renable <= 0;
        _stream_matmul_33_source_21_source_fifo_deq <= 0;
      end 
      _stream_matmul_33_source_21_idle <= _stream_matmul_33_source_21_idle;
      if(_stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_22_source_ram_renable <= 0;
        _stream_matmul_33_source_22_source_fifo_deq <= 0;
      end 
      _stream_matmul_33_source_22_idle <= _stream_matmul_33_source_22_idle;
      if(_stream_matmul_33_stream_oready) begin
        _stream_matmul_33_sink_33_sink_wenable <= 0;
        _stream_matmul_33_sink_33_sink_fifo_enq <= 0;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _stream_matmul_33_sink_34_sink_wenable <= 0;
        _stream_matmul_33_sink_34_sink_fifo_enq <= 0;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_1 <= _stream_matmul_33_stream_ivalid;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_2 <= __stream_matmul_33_stream_ivalid_1;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_3 <= __stream_matmul_33_stream_ivalid_2;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_4 <= __stream_matmul_33_stream_ivalid_3;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_5 <= __stream_matmul_33_stream_ivalid_4;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_6 <= __stream_matmul_33_stream_ivalid_5;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_7 <= __stream_matmul_33_stream_ivalid_6;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_8 <= __stream_matmul_33_stream_ivalid_7;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_9 <= __stream_matmul_33_stream_ivalid_8;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_10 <= __stream_matmul_33_stream_ivalid_9;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_11 <= __stream_matmul_33_stream_ivalid_10;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_12 <= __stream_matmul_33_stream_ivalid_11;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_13 <= __stream_matmul_33_stream_ivalid_12;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_14 <= __stream_matmul_33_stream_ivalid_13;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_15 <= __stream_matmul_33_stream_ivalid_14;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_16 <= __stream_matmul_33_stream_ivalid_15;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_17 <= __stream_matmul_33_stream_ivalid_16;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_18 <= __stream_matmul_33_stream_ivalid_17;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_19 <= __stream_matmul_33_stream_ivalid_18;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_20 <= __stream_matmul_33_stream_ivalid_19;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_21 <= __stream_matmul_33_stream_ivalid_20;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_22 <= __stream_matmul_33_stream_ivalid_21;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_23 <= __stream_matmul_33_stream_ivalid_22;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_24 <= __stream_matmul_33_stream_ivalid_23;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_25 <= __stream_matmul_33_stream_ivalid_24;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_26 <= __stream_matmul_33_stream_ivalid_25;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_27 <= __stream_matmul_33_stream_ivalid_26;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_28 <= __stream_matmul_33_stream_ivalid_27;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_29 <= __stream_matmul_33_stream_ivalid_28;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __stream_matmul_33_stream_ivalid_30 <= __stream_matmul_33_stream_ivalid_29;
      end 
      if(_stream_matmul_33_stream_ivalid && _stream_matmul_33_stream_oready && _counter_reset_cond_1058) begin
        _counter_data_1058 <= 1'sd0;
      end 
      if(_stream_matmul_33_stream_ivalid && _stream_matmul_33_stream_oready) begin
        _counter_data_1058 <= _counter_current_count_1058;
      end 
      if(_stream_matmul_33_stream_ivalid && _stream_matmul_33_stream_oready) begin
        _counter_count_1058 <= (_counter_current_count_1058 >= stream_matmul_33_parameter_0_data - 2'sd1)? _counter_current_count_1058 + 2'sd1 - stream_matmul_33_parameter_0_data : _counter_current_count_1058 + 2'sd1;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _minus_data_1063 <= stream_matmul_33_parameter_0_data - 2'sd1;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _minus_data_1069 <= stream_matmul_33_parameter_0_data - 2'sd1;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _eq_data_1138 <= stream_matmul_33_parameter_1_data == 1'sd0;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _eq_data_1142 <= stream_matmul_33_parameter_2_data == 1'sd0;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _plus_data_1189 <= _cond_data_1107 + stream_matmul_33_parameter_16_data;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _plus_data_1194 <= _cond_data_1107 + stream_matmul_33_parameter_16_data;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _plus_data_1199 <= _cond_data_1119 + stream_matmul_33_parameter_17_data;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _plus_data_1204 <= _cond_data_1131 + stream_matmul_33_parameter_18_data;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _plus_data_1210 <= _cond_data_1108 + stream_matmul_33_parameter_16_data;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _plus_data_1215 <= _cond_data_1108 + stream_matmul_33_parameter_16_data;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _plus_data_1231 <= _cond_data_1120 + stream_matmul_33_parameter_17_data;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _plus_data_1250 <= _cond_data_1132 + stream_matmul_33_parameter_18_data;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1501_pointer_1061 <= _pointer_data_1061;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1503__variable_1137 <= stream_matmul_33_source_20_data;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1506_pointer_1184 <= _pointer_data_1184;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1509_reinterpretcast_1163 <= _reinterpretcast_data_1163;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1514_pointer_1067 <= _pointer_data_1067;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1518_reinterpretcast_1167 <= _reinterpretcast_data_1167;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1523__variable_1057 <= stream_matmul_33__reduce_reset_data;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1550__variable_1052 <= stream_matmul_33_parameter_0_data;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1564_reinterpretcast_1175 <= _reinterpretcast_data_1175;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1569_reinterpretcast_1179 <= _reinterpretcast_data_1179;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1587_cond_1084 <= _cond_data_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1607_cond_1096 <= _cond_data_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1648_cond_1083 <= _cond_data_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1668_cond_1095 <= _cond_data_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _eq_data_1065 <= _counter_data_1058 == _minus_data_1063;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _eq_data_1071 <= _counter_data_1058 == _minus_data_1069;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1502__delay_1501_pointer_1061 <= __delay_data_1501_pointer_1061;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1504_reinterpretcast_1149 <= _reinterpretcast_data_1149;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1507__delay_1506_pointer_1184 <= __delay_data_1506_pointer_1184;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1510__delay_1509_reinterpretcast_1163 <= __delay_data_1509_reinterpretcast_1163;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1512_plus_1189 <= _plus_data_1189;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1515__delay_1514_pointer_1067 <= __delay_data_1514_pointer_1067;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1516_reinterpretcast_1153 <= _reinterpretcast_data_1153;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1519__delay_1518_reinterpretcast_1167 <= __delay_data_1518_reinterpretcast_1167;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1521_plus_1194 <= _plus_data_1194;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1524__delay_1523__variable_1057 <= __delay_data_1523__variable_1057;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1537_plus_1199 <= _plus_data_1199;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1551__delay_1550__variable_1052 <= __delay_data_1550__variable_1052;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1565__delay_1564_reinterpretcast_1175 <= __delay_data_1564_reinterpretcast_1175;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1567_plus_1210 <= _plus_data_1210;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1570__delay_1569_reinterpretcast_1179 <= __delay_data_1569_reinterpretcast_1179;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1572_plus_1215 <= _plus_data_1215;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1574_plus_1231 <= _plus_data_1231;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1588__delay_1587_cond_1084 <= __delay_data_1587_cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1608__delay_1607_cond_1096 <= __delay_data_1607_cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1628_plus_1250 <= _plus_data_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1649__delay_1648_cond_1083 <= __delay_data_1648_cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1669__delay_1668_cond_1095 <= __delay_data_1668_cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1689_plus_1204 <= _plus_data_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _land_data_1066 <= __delay_data_1502__delay_1501_pointer_1061 && _eq_data_1065;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _land_data_1072 <= __delay_data_1515__delay_1514_pointer_1067 && _eq_data_1071;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1505__delay_1504_reinterpretcast_1149 <= __delay_data_1504_reinterpretcast_1149;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1508__delay_1507__delay_1506_pointer_1184 <= __delay_data_1507__delay_1506_pointer_1184;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1511__delay_1510__delay_1509_reinterpretcast_1163 <= __delay_data_1510__delay_1509_reinterpretcast_1163;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1513__delay_1512_plus_1189 <= __delay_data_1512_plus_1189;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1517__delay_1516_reinterpretcast_1153 <= __delay_data_1516_reinterpretcast_1153;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1520__delay_1519__delay_1518_reinterpretcast_1167 <= __delay_data_1519__delay_1518_reinterpretcast_1167;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1522__delay_1521_plus_1194 <= __delay_data_1521_plus_1194;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1525__delay_1524__delay_1523__variable_1057 <= __delay_data_1524__delay_1523__variable_1057;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1538__delay_1537_plus_1199 <= __delay_data_1537_plus_1199;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1552__delay_1551__delay_1550__variable_1052 <= __delay_data_1551__delay_1550__variable_1052;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1566__delay_1565__delay_1564_reinterpretcast_1175 <= __delay_data_1565__delay_1564_reinterpretcast_1175;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1568__delay_1567_plus_1210 <= __delay_data_1567_plus_1210;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1571__delay_1570__delay_1569_reinterpretcast_1179 <= __delay_data_1570__delay_1569_reinterpretcast_1179;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1573__delay_1572_plus_1215 <= __delay_data_1572_plus_1215;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1575__delay_1574_plus_1231 <= __delay_data_1574_plus_1231;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1589__delay_1588__delay_1587_cond_1084 <= __delay_data_1588__delay_1587_cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1609__delay_1608__delay_1607_cond_1096 <= __delay_data_1608__delay_1607_cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1629__delay_1628_plus_1250 <= __delay_data_1628_plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1650__delay_1649__delay_1648_cond_1083 <= __delay_data_1649__delay_1648_cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1670__delay_1669__delay_1668_cond_1095 <= __delay_data_1669__delay_1668_cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1690__delay_1689_plus_1204 <= __delay_data_1689_plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1526__delay_1525__delay_1524____variable_1057 <= __delay_data_1525__delay_1524__delay_1523__variable_1057;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1539__delay_1538__delay_1537_plus_1199 <= __delay_data_1538__delay_1537_plus_1199;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1553__delay_1552__delay_1551____variable_1052 <= __delay_data_1552__delay_1551__delay_1550__variable_1052;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1576__delay_1575__delay_1574_plus_1231 <= __delay_data_1575__delay_1574_plus_1231;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1590__delay_1589__delay_1588___cond_1084 <= __delay_data_1589__delay_1588__delay_1587_cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1610__delay_1609__delay_1608___cond_1096 <= __delay_data_1609__delay_1608__delay_1607_cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1630__delay_1629__delay_1628_plus_1250 <= __delay_data_1629__delay_1628_plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1651__delay_1650__delay_1649___cond_1083 <= __delay_data_1650__delay_1649__delay_1648_cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1671__delay_1670__delay_1669___cond_1095 <= __delay_data_1670__delay_1669__delay_1668_cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1691__delay_1690__delay_1689_plus_1204 <= __delay_data_1690__delay_1689_plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1527__delay_1526__delay_1525____variable_1057 <= __delay_data_1526__delay_1525__delay_1524____variable_1057;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1540__delay_1539__delay_1538___plus_1199 <= __delay_data_1539__delay_1538__delay_1537_plus_1199;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1554__delay_1553__delay_1552____variable_1052 <= __delay_data_1553__delay_1552__delay_1551____variable_1052;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1577__delay_1576__delay_1575___plus_1231 <= __delay_data_1576__delay_1575__delay_1574_plus_1231;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1591__delay_1590__delay_1589___cond_1084 <= __delay_data_1590__delay_1589__delay_1588___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1611__delay_1610__delay_1609___cond_1096 <= __delay_data_1610__delay_1609__delay_1608___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1631__delay_1630__delay_1629___plus_1250 <= __delay_data_1630__delay_1629__delay_1628_plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1652__delay_1651__delay_1650___cond_1083 <= __delay_data_1651__delay_1650__delay_1649___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1672__delay_1671__delay_1670___cond_1095 <= __delay_data_1671__delay_1670__delay_1669___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1692__delay_1691__delay_1690___plus_1204 <= __delay_data_1691__delay_1690__delay_1689_plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1528__delay_1527__delay_1526____variable_1057 <= __delay_data_1527__delay_1526__delay_1525____variable_1057;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1541__delay_1540__delay_1539___plus_1199 <= __delay_data_1540__delay_1539__delay_1538___plus_1199;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1555__delay_1554__delay_1553____variable_1052 <= __delay_data_1554__delay_1553__delay_1552____variable_1052;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1578__delay_1577__delay_1576___plus_1231 <= __delay_data_1577__delay_1576__delay_1575___plus_1231;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1592__delay_1591__delay_1590___cond_1084 <= __delay_data_1591__delay_1590__delay_1589___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1612__delay_1611__delay_1610___cond_1096 <= __delay_data_1611__delay_1610__delay_1609___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1632__delay_1631__delay_1630___plus_1250 <= __delay_data_1631__delay_1630__delay_1629___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1653__delay_1652__delay_1651___cond_1083 <= __delay_data_1652__delay_1651__delay_1650___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1673__delay_1672__delay_1671___cond_1095 <= __delay_data_1672__delay_1671__delay_1670___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1693__delay_1692__delay_1691___plus_1204 <= __delay_data_1692__delay_1691__delay_1690___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1529__delay_1528__delay_1527____variable_1057 <= __delay_data_1528__delay_1527__delay_1526____variable_1057;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1542__delay_1541__delay_1540___plus_1199 <= __delay_data_1541__delay_1540__delay_1539___plus_1199;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1556__delay_1555__delay_1554____variable_1052 <= __delay_data_1555__delay_1554__delay_1553____variable_1052;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1579__delay_1578__delay_1577___plus_1231 <= __delay_data_1578__delay_1577__delay_1576___plus_1231;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1593__delay_1592__delay_1591___cond_1084 <= __delay_data_1592__delay_1591__delay_1590___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1613__delay_1612__delay_1611___cond_1096 <= __delay_data_1612__delay_1611__delay_1610___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1633__delay_1632__delay_1631___plus_1250 <= __delay_data_1632__delay_1631__delay_1630___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1654__delay_1653__delay_1652___cond_1083 <= __delay_data_1653__delay_1652__delay_1651___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1674__delay_1673__delay_1672___cond_1095 <= __delay_data_1673__delay_1672__delay_1671___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1694__delay_1693__delay_1692___plus_1204 <= __delay_data_1693__delay_1692__delay_1691___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1530__delay_1529__delay_1528____variable_1057 <= __delay_data_1529__delay_1528__delay_1527____variable_1057;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1543__delay_1542__delay_1541___plus_1199 <= __delay_data_1542__delay_1541__delay_1540___plus_1199;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1557__delay_1556__delay_1555____variable_1052 <= __delay_data_1556__delay_1555__delay_1554____variable_1052;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1580__delay_1579__delay_1578___plus_1231 <= __delay_data_1579__delay_1578__delay_1577___plus_1231;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1594__delay_1593__delay_1592___cond_1084 <= __delay_data_1593__delay_1592__delay_1591___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1614__delay_1613__delay_1612___cond_1096 <= __delay_data_1613__delay_1612__delay_1611___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1634__delay_1633__delay_1632___plus_1250 <= __delay_data_1633__delay_1632__delay_1631___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1655__delay_1654__delay_1653___cond_1083 <= __delay_data_1654__delay_1653__delay_1652___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1675__delay_1674__delay_1673___cond_1095 <= __delay_data_1674__delay_1673__delay_1672___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1695__delay_1694__delay_1693___plus_1204 <= __delay_data_1694__delay_1693__delay_1692___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1531__delay_1530__delay_1529____variable_1057 <= __delay_data_1530__delay_1529__delay_1528____variable_1057;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1544__delay_1543__delay_1542___plus_1199 <= __delay_data_1543__delay_1542__delay_1541___plus_1199;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1558__delay_1557__delay_1556____variable_1052 <= __delay_data_1557__delay_1556__delay_1555____variable_1052;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1581__delay_1580__delay_1579___plus_1231 <= __delay_data_1580__delay_1579__delay_1578___plus_1231;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1595__delay_1594__delay_1593___cond_1084 <= __delay_data_1594__delay_1593__delay_1592___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1615__delay_1614__delay_1613___cond_1096 <= __delay_data_1614__delay_1613__delay_1612___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1635__delay_1634__delay_1633___plus_1250 <= __delay_data_1634__delay_1633__delay_1632___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1656__delay_1655__delay_1654___cond_1083 <= __delay_data_1655__delay_1654__delay_1653___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1676__delay_1675__delay_1674___cond_1095 <= __delay_data_1675__delay_1674__delay_1673___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1696__delay_1695__delay_1694___plus_1204 <= __delay_data_1695__delay_1694__delay_1693___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1532__delay_1531__delay_1530____variable_1057 <= __delay_data_1531__delay_1530__delay_1529____variable_1057;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1545__delay_1544__delay_1543___plus_1199 <= __delay_data_1544__delay_1543__delay_1542___plus_1199;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1559__delay_1558__delay_1557____variable_1052 <= __delay_data_1558__delay_1557__delay_1556____variable_1052;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1582__delay_1581__delay_1580___plus_1231 <= __delay_data_1581__delay_1580__delay_1579___plus_1231;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1596__delay_1595__delay_1594___cond_1084 <= __delay_data_1595__delay_1594__delay_1593___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1616__delay_1615__delay_1614___cond_1096 <= __delay_data_1615__delay_1614__delay_1613___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1636__delay_1635__delay_1634___plus_1250 <= __delay_data_1635__delay_1634__delay_1633___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1657__delay_1656__delay_1655___cond_1083 <= __delay_data_1656__delay_1655__delay_1654___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1677__delay_1676__delay_1675___cond_1095 <= __delay_data_1676__delay_1675__delay_1674___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1697__delay_1696__delay_1695___plus_1204 <= __delay_data_1696__delay_1695__delay_1694___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1533__delay_1532__delay_1531____variable_1057 <= __delay_data_1532__delay_1531__delay_1530____variable_1057;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1546__delay_1545__delay_1544___plus_1199 <= __delay_data_1545__delay_1544__delay_1543___plus_1199;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1560__delay_1559__delay_1558____variable_1052 <= __delay_data_1559__delay_1558__delay_1557____variable_1052;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1583__delay_1582__delay_1581___plus_1231 <= __delay_data_1582__delay_1581__delay_1580___plus_1231;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1597__delay_1596__delay_1595___cond_1084 <= __delay_data_1596__delay_1595__delay_1594___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1617__delay_1616__delay_1615___cond_1096 <= __delay_data_1616__delay_1615__delay_1614___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1637__delay_1636__delay_1635___plus_1250 <= __delay_data_1636__delay_1635__delay_1634___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1658__delay_1657__delay_1656___cond_1083 <= __delay_data_1657__delay_1656__delay_1655___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1678__delay_1677__delay_1676___cond_1095 <= __delay_data_1677__delay_1676__delay_1675___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1698__delay_1697__delay_1696___plus_1204 <= __delay_data_1697__delay_1696__delay_1695___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1534__delay_1533__delay_1532____variable_1057 <= __delay_data_1533__delay_1532__delay_1531____variable_1057;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1547__delay_1546__delay_1545___plus_1199 <= __delay_data_1546__delay_1545__delay_1544___plus_1199;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1561__delay_1560__delay_1559____variable_1052 <= __delay_data_1560__delay_1559__delay_1558____variable_1052;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1584__delay_1583__delay_1582___plus_1231 <= __delay_data_1583__delay_1582__delay_1581___plus_1231;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1598__delay_1597__delay_1596___cond_1084 <= __delay_data_1597__delay_1596__delay_1595___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1618__delay_1617__delay_1616___cond_1096 <= __delay_data_1617__delay_1616__delay_1615___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1638__delay_1637__delay_1636___plus_1250 <= __delay_data_1637__delay_1636__delay_1635___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1659__delay_1658__delay_1657___cond_1083 <= __delay_data_1658__delay_1657__delay_1656___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1679__delay_1678__delay_1677___cond_1095 <= __delay_data_1678__delay_1677__delay_1676___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1699__delay_1698__delay_1697___plus_1204 <= __delay_data_1698__delay_1697__delay_1696___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1535__delay_1534__delay_1533____variable_1057 <= __delay_data_1534__delay_1533__delay_1532____variable_1057;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1548__delay_1547__delay_1546___plus_1199 <= __delay_data_1547__delay_1546__delay_1545___plus_1199;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1562__delay_1561__delay_1560____variable_1052 <= __delay_data_1561__delay_1560__delay_1559____variable_1052;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1585__delay_1584__delay_1583___plus_1231 <= __delay_data_1584__delay_1583__delay_1582___plus_1231;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1599__delay_1598__delay_1597___cond_1084 <= __delay_data_1598__delay_1597__delay_1596___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1619__delay_1618__delay_1617___cond_1096 <= __delay_data_1618__delay_1617__delay_1616___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1639__delay_1638__delay_1637___plus_1250 <= __delay_data_1638__delay_1637__delay_1636___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1660__delay_1659__delay_1658___cond_1083 <= __delay_data_1659__delay_1658__delay_1657___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1680__delay_1679__delay_1678___cond_1095 <= __delay_data_1679__delay_1678__delay_1677___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1700__delay_1699__delay_1698___plus_1204 <= __delay_data_1699__delay_1698__delay_1697___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1536__delay_1535__delay_1534____variable_1057 <= __delay_data_1535__delay_1534__delay_1533____variable_1057;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1549__delay_1548__delay_1547___plus_1199 <= __delay_data_1548__delay_1547__delay_1546___plus_1199;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1563__delay_1562__delay_1561____variable_1052 <= __delay_data_1562__delay_1561__delay_1560____variable_1052;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1586__delay_1585__delay_1584___plus_1231 <= __delay_data_1585__delay_1584__delay_1583___plus_1231;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1600__delay_1599__delay_1598___cond_1084 <= __delay_data_1599__delay_1598__delay_1597___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1620__delay_1619__delay_1618___cond_1096 <= __delay_data_1619__delay_1618__delay_1617___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1640__delay_1639__delay_1638___plus_1250 <= __delay_data_1639__delay_1638__delay_1637___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1661__delay_1660__delay_1659___cond_1083 <= __delay_data_1660__delay_1659__delay_1658___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1681__delay_1680__delay_1679___cond_1095 <= __delay_data_1680__delay_1679__delay_1678___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1701__delay_1700__delay_1699___plus_1204 <= __delay_data_1700__delay_1699__delay_1698___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1601__delay_1600__delay_1599___cond_1084 <= __delay_data_1600__delay_1599__delay_1598___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1621__delay_1620__delay_1619___cond_1096 <= __delay_data_1620__delay_1619__delay_1618___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1641__delay_1640__delay_1639___plus_1250 <= __delay_data_1640__delay_1639__delay_1638___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1662__delay_1661__delay_1660___cond_1083 <= __delay_data_1661__delay_1660__delay_1659___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1682__delay_1681__delay_1680___cond_1095 <= __delay_data_1681__delay_1680__delay_1679___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1702__delay_1701__delay_1700___plus_1204 <= __delay_data_1701__delay_1700__delay_1699___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1602__delay_1601__delay_1600___cond_1084 <= __delay_data_1601__delay_1600__delay_1599___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1622__delay_1621__delay_1620___cond_1096 <= __delay_data_1621__delay_1620__delay_1619___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1642__delay_1641__delay_1640___plus_1250 <= __delay_data_1641__delay_1640__delay_1639___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1663__delay_1662__delay_1661___cond_1083 <= __delay_data_1662__delay_1661__delay_1660___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1683__delay_1682__delay_1681___cond_1095 <= __delay_data_1682__delay_1681__delay_1680___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1703__delay_1702__delay_1701___plus_1204 <= __delay_data_1702__delay_1701__delay_1700___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1603__delay_1602__delay_1601___cond_1084 <= __delay_data_1602__delay_1601__delay_1600___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1623__delay_1622__delay_1621___cond_1096 <= __delay_data_1622__delay_1621__delay_1620___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1643__delay_1642__delay_1641___plus_1250 <= __delay_data_1642__delay_1641__delay_1640___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1664__delay_1663__delay_1662___cond_1083 <= __delay_data_1663__delay_1662__delay_1661___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1684__delay_1683__delay_1682___cond_1095 <= __delay_data_1683__delay_1682__delay_1681___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1704__delay_1703__delay_1702___plus_1204 <= __delay_data_1703__delay_1702__delay_1701___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1604__delay_1603__delay_1602___cond_1084 <= __delay_data_1603__delay_1602__delay_1601___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1624__delay_1623__delay_1622___cond_1096 <= __delay_data_1623__delay_1622__delay_1621___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1644__delay_1643__delay_1642___plus_1250 <= __delay_data_1643__delay_1642__delay_1641___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1665__delay_1664__delay_1663___cond_1083 <= __delay_data_1664__delay_1663__delay_1662___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1685__delay_1684__delay_1683___cond_1095 <= __delay_data_1684__delay_1683__delay_1682___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1705__delay_1704__delay_1703___plus_1204 <= __delay_data_1704__delay_1703__delay_1702___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1605__delay_1604__delay_1603___cond_1084 <= __delay_data_1604__delay_1603__delay_1602___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1625__delay_1624__delay_1623___cond_1096 <= __delay_data_1624__delay_1623__delay_1622___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1645__delay_1644__delay_1643___plus_1250 <= __delay_data_1644__delay_1643__delay_1642___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1666__delay_1665__delay_1664___cond_1083 <= __delay_data_1665__delay_1664__delay_1663___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1686__delay_1685__delay_1684___cond_1095 <= __delay_data_1685__delay_1684__delay_1683___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1706__delay_1705__delay_1704___plus_1204 <= __delay_data_1705__delay_1704__delay_1703___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1606__delay_1605__delay_1604___cond_1084 <= __delay_data_1605__delay_1604__delay_1603___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1626__delay_1625__delay_1624___cond_1096 <= __delay_data_1625__delay_1624__delay_1623___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1646__delay_1645__delay_1644___plus_1250 <= __delay_data_1645__delay_1644__delay_1643___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1667__delay_1666__delay_1665___cond_1083 <= __delay_data_1666__delay_1665__delay_1664___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1687__delay_1686__delay_1685___cond_1095 <= __delay_data_1686__delay_1685__delay_1684___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1707__delay_1706__delay_1705___plus_1204 <= __delay_data_1706__delay_1705__delay_1704___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _plus_data_1202 <= __substreamoutput_data_1200 + __delay_data_1667__delay_1666__delay_1665___cond_1083;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _plus_data_1234 <= __substreamoutput_data_1232 + __delay_data_1606__delay_1605__delay_1604___cond_1084;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1627__delay_1626__delay_1625___cond_1096 <= __delay_data_1626__delay_1625__delay_1624___cond_1096;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1647__delay_1646__delay_1645___plus_1250 <= __delay_data_1646__delay_1645__delay_1644___plus_1250;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1688__delay_1687__delay_1686___cond_1095 <= __delay_data_1687__delay_1686__delay_1685___cond_1095;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1708__delay_1707__delay_1706___plus_1204 <= __delay_data_1707__delay_1706__delay_1705___plus_1204;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1709__substreamoutput_1201 <= __substreamoutput_data_1201;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1710__delay_1709__substreamoutput_1201 <= __delay_data_1709__substreamoutput_1201;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1711__delay_1710____substreamoutput_1201 <= __delay_data_1710__delay_1709__substreamoutput_1201;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1712__delay_1711____substreamoutput_1201 <= __delay_data_1711__delay_1710____substreamoutput_1201;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1713__delay_1712____substreamoutput_1201 <= __delay_data_1712__delay_1711____substreamoutput_1201;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1714__delay_1713____substreamoutput_1201 <= __delay_data_1713__delay_1712____substreamoutput_1201;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1715__delay_1714____substreamoutput_1201 <= __delay_data_1714__delay_1713____substreamoutput_1201;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1716__delay_1715____substreamoutput_1201 <= __delay_data_1715__delay_1714____substreamoutput_1201;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1717__delay_1716____substreamoutput_1201 <= __delay_data_1716__delay_1715____substreamoutput_1201;
      end 
      if(_stream_matmul_33_stream_oready) begin
        __delay_data_1718__delay_1717____substreamoutput_1201 <= __delay_data_1717__delay_1716____substreamoutput_1201;
      end 
      if(_set_flag_1670) begin
        _stream_matmul_33_parameter_0_next_parameter_data <= cparam_matmul_33_stream_reduce_size;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1052 <= _stream_matmul_33_parameter_0_next_parameter_data;
      end 
      if(_set_flag_1671) begin
        _stream_matmul_33_parameter_1_next_parameter_data <= matmul_33_col_select;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1053 <= _stream_matmul_33_parameter_1_next_parameter_data;
      end 
      if(_set_flag_1672) begin
        _stream_matmul_33_parameter_2_next_parameter_data <= matmul_33_row_select_buf;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1054 <= _stream_matmul_33_parameter_2_next_parameter_data;
      end 
      if(_set_flag_1673) begin
        _stream_matmul_33_parameter_3_next_parameter_data <= matmul_33_stream_pad_masks;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1055 <= _stream_matmul_33_parameter_3_next_parameter_data;
      end 
      if(_set_flag_1674) begin
        _stream_matmul_33_parameter_4_next_parameter_data <= cparam_matmul_33_stream_omit_mask;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1056 <= _stream_matmul_33_parameter_4_next_parameter_data;
      end 
      if(_set_flag_1675) begin
        _stream_matmul_33_parameter_6_next_parameter_data <= cparam_matmul_33_bias_scala;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1073 <= _stream_matmul_33_parameter_6_next_parameter_data;
      end 
      if(_set_flag_1676) begin
        _stream_matmul_33_source_7_source_mode <= 5'b10;
        _stream_matmul_33_source_7_source_offset <= (cparam_matmul_33_bias_num == 1)? 0 : matmul_33_och_count_buf;
      end 
      if(_set_flag_1676) begin
        _source_stream_matmul_33_source_7_pat_size_0 <= cparam_matmul_33_stream_reduce_size;
        _source_stream_matmul_33_source_7_pat_stride_0 <= 0;
      end 
      if(_set_flag_1676) begin
        _source_stream_matmul_33_source_7_pat_size_1 <= matmul_33_next_stream_num_ops;
        _source_stream_matmul_33_source_7_pat_stride_1 <= (cparam_matmul_33_bias_num == 1)? 0 : 1;
      end 
      if(_set_flag_1676) begin
        _source_stream_matmul_33_source_7_pat_size_2 <= 1;
        _source_stream_matmul_33_source_7_pat_stride_2 <= 0;
      end 
      if(_set_flag_1676) begin
        _source_stream_matmul_33_source_7_pat_size_3 <= 1;
        _source_stream_matmul_33_source_7_pat_stride_3 <= 0;
      end 
      if(_set_flag_1676) begin
        _stream_matmul_33_source_7_source_sel <= 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_7_source_offset_buf <= _stream_matmul_33_source_7_source_offset;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_count_0 <= _source_stream_matmul_33_source_7_pat_size_0 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_count_1 <= _source_stream_matmul_33_source_7_pat_size_1 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_count_2 <= _source_stream_matmul_33_source_7_pat_size_2 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_count_3 <= _source_stream_matmul_33_source_7_pat_size_3 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_size_buf_0 <= _source_stream_matmul_33_source_7_pat_size_0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_size_buf_1 <= _source_stream_matmul_33_source_7_pat_size_1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_size_buf_2 <= _source_stream_matmul_33_source_7_pat_size_2;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_size_buf_3 <= _source_stream_matmul_33_source_7_pat_size_3;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_stride_buf_0 <= _source_stream_matmul_33_source_7_pat_stride_0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_stride_buf_1 <= _source_stream_matmul_33_source_7_pat_stride_1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_stride_buf_2 <= _source_stream_matmul_33_source_7_pat_stride_2;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_stride_buf_3 <= _source_stream_matmul_33_source_7_pat_stride_3;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_source_busy && _stream_matmul_33_is_root) begin
        __variable_wdata_1074 <= _stream_matmul_33_source_7_source_ram_rdata;
      end 
      if((_stream_matmul_33_source_7_source_pat_fsm_0 == 1) && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_7_idle <= 0;
        _stream_matmul_33_source_7_source_ram_raddr <= _stream_matmul_33_source_7_source_pat_all_offset;
        _stream_matmul_33_source_7_source_ram_renable <= 1;
      end 
      if((_stream_matmul_33_source_7_source_pat_fsm_0 == 1) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_cur_offset_0 <= _source_stream_matmul_33_source_7_pat_cur_offset_0 + _source_stream_matmul_33_source_7_pat_stride_buf_0;
        _source_stream_matmul_33_source_7_pat_count_0 <= _source_stream_matmul_33_source_7_pat_count_0 - 1;
      end 
      if((_stream_matmul_33_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_33_source_7_pat_count_0 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_cur_offset_0 <= 0;
        _source_stream_matmul_33_source_7_pat_count_0 <= _source_stream_matmul_33_source_7_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_33_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_33_source_7_pat_count_0 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_cur_offset_1 <= _source_stream_matmul_33_source_7_pat_cur_offset_1 + _source_stream_matmul_33_source_7_pat_stride_buf_1;
        _source_stream_matmul_33_source_7_pat_count_1 <= _source_stream_matmul_33_source_7_pat_count_1 - 1;
      end 
      if((_stream_matmul_33_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_33_source_7_pat_count_0 == 0) && (_source_stream_matmul_33_source_7_pat_count_1 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_cur_offset_1 <= 0;
        _source_stream_matmul_33_source_7_pat_count_1 <= _source_stream_matmul_33_source_7_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_33_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_33_source_7_pat_count_0 == 0) && (_source_stream_matmul_33_source_7_pat_count_1 == 0)) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_cur_offset_2 <= _source_stream_matmul_33_source_7_pat_cur_offset_2 + _source_stream_matmul_33_source_7_pat_stride_buf_2;
        _source_stream_matmul_33_source_7_pat_count_2 <= _source_stream_matmul_33_source_7_pat_count_2 - 1;
      end 
      if((_stream_matmul_33_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_33_source_7_pat_count_0 == 0) && (_source_stream_matmul_33_source_7_pat_count_1 == 0)) && (_source_stream_matmul_33_source_7_pat_count_2 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_cur_offset_2 <= 0;
        _source_stream_matmul_33_source_7_pat_count_2 <= _source_stream_matmul_33_source_7_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_33_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_33_source_7_pat_count_0 == 0) && (_source_stream_matmul_33_source_7_pat_count_1 == 0) && (_source_stream_matmul_33_source_7_pat_count_2 == 0)) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_cur_offset_3 <= _source_stream_matmul_33_source_7_pat_cur_offset_3 + _source_stream_matmul_33_source_7_pat_stride_buf_3;
        _source_stream_matmul_33_source_7_pat_count_3 <= _source_stream_matmul_33_source_7_pat_count_3 - 1;
      end 
      if((_stream_matmul_33_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_33_source_7_pat_count_0 == 0) && (_source_stream_matmul_33_source_7_pat_count_1 == 0) && (_source_stream_matmul_33_source_7_pat_count_2 == 0)) && (_source_stream_matmul_33_source_7_pat_count_3 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_7_pat_cur_offset_3 <= 0;
        _source_stream_matmul_33_source_7_pat_count_3 <= _source_stream_matmul_33_source_7_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_33_source_7_source_pat_fsm_0 == 1) && _stream_matmul_33_source_stop && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_7_source_ram_renable <= 0;
        _stream_matmul_33_source_7_idle <= 1;
      end 
      if((_stream_matmul_33_source_7_source_pat_fsm_0 == 2) && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_7_source_ram_renable <= 0;
        _stream_matmul_33_source_7_idle <= 1;
      end 
      if(_set_flag_1679) begin
        _stream_matmul_33_parameter_8_next_parameter_data <= cparam_matmul_33_scale_scala;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1085 <= _stream_matmul_33_parameter_8_next_parameter_data;
      end 
      if(_set_flag_1680) begin
        _stream_matmul_33_source_9_source_mode <= 5'b10;
        _stream_matmul_33_source_9_source_offset <= (cparam_matmul_33_scale_num == 1)? 0 : matmul_33_och_count_buf;
      end 
      if(_set_flag_1680) begin
        _source_stream_matmul_33_source_9_pat_size_0 <= cparam_matmul_33_stream_reduce_size;
        _source_stream_matmul_33_source_9_pat_stride_0 <= 0;
      end 
      if(_set_flag_1680) begin
        _source_stream_matmul_33_source_9_pat_size_1 <= matmul_33_next_stream_num_ops;
        _source_stream_matmul_33_source_9_pat_stride_1 <= (cparam_matmul_33_scale_num == 1)? 0 : 1;
      end 
      if(_set_flag_1680) begin
        _source_stream_matmul_33_source_9_pat_size_2 <= 1;
        _source_stream_matmul_33_source_9_pat_stride_2 <= 0;
      end 
      if(_set_flag_1680) begin
        _source_stream_matmul_33_source_9_pat_size_3 <= 1;
        _source_stream_matmul_33_source_9_pat_stride_3 <= 0;
      end 
      if(_set_flag_1680) begin
        _stream_matmul_33_source_9_source_sel <= 2;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_9_source_offset_buf <= _stream_matmul_33_source_9_source_offset;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_count_0 <= _source_stream_matmul_33_source_9_pat_size_0 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_count_1 <= _source_stream_matmul_33_source_9_pat_size_1 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_count_2 <= _source_stream_matmul_33_source_9_pat_size_2 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_count_3 <= _source_stream_matmul_33_source_9_pat_size_3 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_size_buf_0 <= _source_stream_matmul_33_source_9_pat_size_0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_size_buf_1 <= _source_stream_matmul_33_source_9_pat_size_1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_size_buf_2 <= _source_stream_matmul_33_source_9_pat_size_2;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_size_buf_3 <= _source_stream_matmul_33_source_9_pat_size_3;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_stride_buf_0 <= _source_stream_matmul_33_source_9_pat_stride_0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_stride_buf_1 <= _source_stream_matmul_33_source_9_pat_stride_1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_stride_buf_2 <= _source_stream_matmul_33_source_9_pat_stride_2;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_stride_buf_3 <= _source_stream_matmul_33_source_9_pat_stride_3;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_source_busy && _stream_matmul_33_is_root) begin
        __variable_wdata_1086 <= _stream_matmul_33_source_9_source_ram_rdata;
      end 
      if((_stream_matmul_33_source_9_source_pat_fsm_1 == 1) && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_9_idle <= 0;
        _stream_matmul_33_source_9_source_ram_raddr <= _stream_matmul_33_source_9_source_pat_all_offset;
        _stream_matmul_33_source_9_source_ram_renable <= 1;
      end 
      if((_stream_matmul_33_source_9_source_pat_fsm_1 == 1) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_cur_offset_0 <= _source_stream_matmul_33_source_9_pat_cur_offset_0 + _source_stream_matmul_33_source_9_pat_stride_buf_0;
        _source_stream_matmul_33_source_9_pat_count_0 <= _source_stream_matmul_33_source_9_pat_count_0 - 1;
      end 
      if((_stream_matmul_33_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_33_source_9_pat_count_0 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_cur_offset_0 <= 0;
        _source_stream_matmul_33_source_9_pat_count_0 <= _source_stream_matmul_33_source_9_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_33_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_33_source_9_pat_count_0 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_cur_offset_1 <= _source_stream_matmul_33_source_9_pat_cur_offset_1 + _source_stream_matmul_33_source_9_pat_stride_buf_1;
        _source_stream_matmul_33_source_9_pat_count_1 <= _source_stream_matmul_33_source_9_pat_count_1 - 1;
      end 
      if((_stream_matmul_33_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_33_source_9_pat_count_0 == 0) && (_source_stream_matmul_33_source_9_pat_count_1 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_cur_offset_1 <= 0;
        _source_stream_matmul_33_source_9_pat_count_1 <= _source_stream_matmul_33_source_9_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_33_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_33_source_9_pat_count_0 == 0) && (_source_stream_matmul_33_source_9_pat_count_1 == 0)) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_cur_offset_2 <= _source_stream_matmul_33_source_9_pat_cur_offset_2 + _source_stream_matmul_33_source_9_pat_stride_buf_2;
        _source_stream_matmul_33_source_9_pat_count_2 <= _source_stream_matmul_33_source_9_pat_count_2 - 1;
      end 
      if((_stream_matmul_33_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_33_source_9_pat_count_0 == 0) && (_source_stream_matmul_33_source_9_pat_count_1 == 0)) && (_source_stream_matmul_33_source_9_pat_count_2 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_cur_offset_2 <= 0;
        _source_stream_matmul_33_source_9_pat_count_2 <= _source_stream_matmul_33_source_9_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_33_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_33_source_9_pat_count_0 == 0) && (_source_stream_matmul_33_source_9_pat_count_1 == 0) && (_source_stream_matmul_33_source_9_pat_count_2 == 0)) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_cur_offset_3 <= _source_stream_matmul_33_source_9_pat_cur_offset_3 + _source_stream_matmul_33_source_9_pat_stride_buf_3;
        _source_stream_matmul_33_source_9_pat_count_3 <= _source_stream_matmul_33_source_9_pat_count_3 - 1;
      end 
      if((_stream_matmul_33_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_33_source_9_pat_count_0 == 0) && (_source_stream_matmul_33_source_9_pat_count_1 == 0) && (_source_stream_matmul_33_source_9_pat_count_2 == 0)) && (_source_stream_matmul_33_source_9_pat_count_3 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_9_pat_cur_offset_3 <= 0;
        _source_stream_matmul_33_source_9_pat_count_3 <= _source_stream_matmul_33_source_9_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_33_source_9_source_pat_fsm_1 == 1) && _stream_matmul_33_source_stop && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_9_source_ram_renable <= 0;
        _stream_matmul_33_source_9_idle <= 1;
      end 
      if((_stream_matmul_33_source_9_source_pat_fsm_1 == 2) && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_9_source_ram_renable <= 0;
        _stream_matmul_33_source_9_idle <= 1;
      end 
      if(_set_flag_1683) begin
        _stream_matmul_33_parameter_10_next_parameter_data <= 1;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1097 <= _stream_matmul_33_parameter_10_next_parameter_data;
      end 
      if(_set_flag_1684) begin
        _stream_matmul_33_source_11_source_mode <= 5'b0;
        _stream_matmul_33_source_11_source_empty_data <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_stream_oready && !(|(_stream_matmul_33_source_11_source_mode & 5'b0))) begin
        _stream_matmul_33_source_11_idle <= 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_stream_oready && !(|(_stream_matmul_33_source_11_source_mode & 5'b0)) && _stream_matmul_33_is_root) begin
        __variable_wdata_1098 <= _stream_matmul_33_source_11_source_empty_data;
      end 
      if(_set_flag_1685) begin
        _stream_matmul_33_parameter_12_next_parameter_data <= 1;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1109 <= _stream_matmul_33_parameter_12_next_parameter_data;
      end 
      if(_set_flag_1686) begin
        _stream_matmul_33_source_13_source_mode <= 5'b0;
        _stream_matmul_33_source_13_source_empty_data <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_stream_oready && !(|(_stream_matmul_33_source_13_source_mode & 5'b0))) begin
        _stream_matmul_33_source_13_idle <= 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_stream_oready && !(|(_stream_matmul_33_source_13_source_mode & 5'b0)) && _stream_matmul_33_is_root) begin
        __variable_wdata_1110 <= _stream_matmul_33_source_13_source_empty_data;
      end 
      if(_set_flag_1687) begin
        _stream_matmul_33_parameter_14_next_parameter_data <= 1;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1121 <= _stream_matmul_33_parameter_14_next_parameter_data;
      end 
      if(_set_flag_1688) begin
        _stream_matmul_33_source_15_source_mode <= 5'b0;
        _stream_matmul_33_source_15_source_empty_data <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_stream_oready && !(|(_stream_matmul_33_source_15_source_mode & 5'b0))) begin
        _stream_matmul_33_source_15_idle <= 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_stream_oready && !(|(_stream_matmul_33_source_15_source_mode & 5'b0)) && _stream_matmul_33_is_root) begin
        __variable_wdata_1122 <= _stream_matmul_33_source_15_source_empty_data;
      end 
      if(_set_flag_1689) begin
        _stream_matmul_33_parameter_16_next_parameter_data <= cparam_matmul_33_cshamt_mul_value;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1133 <= _stream_matmul_33_parameter_16_next_parameter_data;
      end 
      if(_set_flag_1690) begin
        _stream_matmul_33_parameter_17_next_parameter_data <= cparam_matmul_33_cshamt_sum_value;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1134 <= _stream_matmul_33_parameter_17_next_parameter_data;
      end 
      if(_set_flag_1691) begin
        _stream_matmul_33_parameter_18_next_parameter_data <= cparam_matmul_33_cshamt_out_value;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1135 <= _stream_matmul_33_parameter_18_next_parameter_data;
      end 
      if(_set_flag_1692) begin
        _stream_matmul_33_parameter_19_next_parameter_data <= cparam_matmul_33_act_func_index;
      end 
      if(_stream_matmul_33_source_start) begin
        __variable_wdata_1136 <= _stream_matmul_33_parameter_19_next_parameter_data;
      end 
      if(_set_flag_1693) begin
        _stream_matmul_33_source_20_source_mode <= 5'b10;
        _stream_matmul_33_source_20_source_offset <= matmul_33_stream_act_local_0 + matmul_33_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_1693) begin
        _source_stream_matmul_33_source_20_pat_size_0 <= cparam_matmul_33_stream_reduce_size;
        _source_stream_matmul_33_source_20_pat_stride_0 <= 1;
      end 
      if(_set_flag_1693) begin
        _source_stream_matmul_33_source_20_pat_size_1 <= matmul_33_next_stream_num_ops;
        _source_stream_matmul_33_source_20_pat_stride_1 <= 0;
      end 
      if(_set_flag_1693) begin
        _source_stream_matmul_33_source_20_pat_size_2 <= 1;
        _source_stream_matmul_33_source_20_pat_stride_2 <= 0;
      end 
      if(_set_flag_1693) begin
        _source_stream_matmul_33_source_20_pat_size_3 <= 1;
        _source_stream_matmul_33_source_20_pat_stride_3 <= 0;
      end 
      if(_set_flag_1693) begin
        _stream_matmul_33_source_20_source_sel <= 3;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_20_source_offset_buf <= _stream_matmul_33_source_20_source_offset;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_count_0 <= _source_stream_matmul_33_source_20_pat_size_0 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_count_1 <= _source_stream_matmul_33_source_20_pat_size_1 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_count_2 <= _source_stream_matmul_33_source_20_pat_size_2 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_count_3 <= _source_stream_matmul_33_source_20_pat_size_3 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_size_buf_0 <= _source_stream_matmul_33_source_20_pat_size_0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_size_buf_1 <= _source_stream_matmul_33_source_20_pat_size_1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_size_buf_2 <= _source_stream_matmul_33_source_20_pat_size_2;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_size_buf_3 <= _source_stream_matmul_33_source_20_pat_size_3;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_stride_buf_0 <= _source_stream_matmul_33_source_20_pat_stride_0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_stride_buf_1 <= _source_stream_matmul_33_source_20_pat_stride_1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_stride_buf_2 <= _source_stream_matmul_33_source_20_pat_stride_2;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_stride_buf_3 <= _source_stream_matmul_33_source_20_pat_stride_3;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_source_busy && _stream_matmul_33_is_root) begin
        __variable_wdata_1137 <= _stream_matmul_33_source_20_source_ram_rdata;
      end 
      if((_stream_matmul_33_source_20_source_pat_fsm_2 == 1) && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_20_idle <= 0;
        _stream_matmul_33_source_20_source_ram_raddr <= _stream_matmul_33_source_20_source_pat_all_offset;
        _stream_matmul_33_source_20_source_ram_renable <= 1;
      end 
      if((_stream_matmul_33_source_20_source_pat_fsm_2 == 1) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_cur_offset_0 <= _source_stream_matmul_33_source_20_pat_cur_offset_0 + _source_stream_matmul_33_source_20_pat_stride_buf_0;
        _source_stream_matmul_33_source_20_pat_count_0 <= _source_stream_matmul_33_source_20_pat_count_0 - 1;
      end 
      if((_stream_matmul_33_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_33_source_20_pat_count_0 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_cur_offset_0 <= 0;
        _source_stream_matmul_33_source_20_pat_count_0 <= _source_stream_matmul_33_source_20_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_33_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_33_source_20_pat_count_0 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_cur_offset_1 <= _source_stream_matmul_33_source_20_pat_cur_offset_1 + _source_stream_matmul_33_source_20_pat_stride_buf_1;
        _source_stream_matmul_33_source_20_pat_count_1 <= _source_stream_matmul_33_source_20_pat_count_1 - 1;
      end 
      if((_stream_matmul_33_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_33_source_20_pat_count_0 == 0) && (_source_stream_matmul_33_source_20_pat_count_1 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_cur_offset_1 <= 0;
        _source_stream_matmul_33_source_20_pat_count_1 <= _source_stream_matmul_33_source_20_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_33_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_33_source_20_pat_count_0 == 0) && (_source_stream_matmul_33_source_20_pat_count_1 == 0)) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_cur_offset_2 <= _source_stream_matmul_33_source_20_pat_cur_offset_2 + _source_stream_matmul_33_source_20_pat_stride_buf_2;
        _source_stream_matmul_33_source_20_pat_count_2 <= _source_stream_matmul_33_source_20_pat_count_2 - 1;
      end 
      if((_stream_matmul_33_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_33_source_20_pat_count_0 == 0) && (_source_stream_matmul_33_source_20_pat_count_1 == 0)) && (_source_stream_matmul_33_source_20_pat_count_2 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_cur_offset_2 <= 0;
        _source_stream_matmul_33_source_20_pat_count_2 <= _source_stream_matmul_33_source_20_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_33_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_33_source_20_pat_count_0 == 0) && (_source_stream_matmul_33_source_20_pat_count_1 == 0) && (_source_stream_matmul_33_source_20_pat_count_2 == 0)) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_cur_offset_3 <= _source_stream_matmul_33_source_20_pat_cur_offset_3 + _source_stream_matmul_33_source_20_pat_stride_buf_3;
        _source_stream_matmul_33_source_20_pat_count_3 <= _source_stream_matmul_33_source_20_pat_count_3 - 1;
      end 
      if((_stream_matmul_33_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_33_source_20_pat_count_0 == 0) && (_source_stream_matmul_33_source_20_pat_count_1 == 0) && (_source_stream_matmul_33_source_20_pat_count_2 == 0)) && (_source_stream_matmul_33_source_20_pat_count_3 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_20_pat_cur_offset_3 <= 0;
        _source_stream_matmul_33_source_20_pat_count_3 <= _source_stream_matmul_33_source_20_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_33_source_20_source_pat_fsm_2 == 1) && _stream_matmul_33_source_stop && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_20_source_ram_renable <= 0;
        _stream_matmul_33_source_20_idle <= 1;
      end 
      if((_stream_matmul_33_source_20_source_pat_fsm_2 == 2) && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_20_source_ram_renable <= 0;
        _stream_matmul_33_source_20_idle <= 1;
      end 
      if(_set_flag_1696) begin
        _stream_matmul_33_source_21_source_mode <= 5'b10;
        _stream_matmul_33_source_21_source_offset <= matmul_33_filter_page_comp_offset_buf;
      end 
      if(_set_flag_1696) begin
        _source_stream_matmul_33_source_21_pat_size_0 <= cparam_matmul_33_stream_reduce_size;
        _source_stream_matmul_33_source_21_pat_stride_0 <= 1;
      end 
      if(_set_flag_1696) begin
        _source_stream_matmul_33_source_21_pat_size_1 <= matmul_33_next_stream_num_ops;
        _source_stream_matmul_33_source_21_pat_stride_1 <= cparam_matmul_33_stream_aligned_reduce_size;
      end 
      if(_set_flag_1696) begin
        _source_stream_matmul_33_source_21_pat_size_2 <= 1;
        _source_stream_matmul_33_source_21_pat_stride_2 <= 0;
      end 
      if(_set_flag_1696) begin
        _source_stream_matmul_33_source_21_pat_size_3 <= 1;
        _source_stream_matmul_33_source_21_pat_stride_3 <= 0;
      end 
      if(_set_flag_1696) begin
        _stream_matmul_33_source_21_source_sel <= 4;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_21_source_offset_buf <= _stream_matmul_33_source_21_source_offset;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_count_0 <= _source_stream_matmul_33_source_21_pat_size_0 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_count_1 <= _source_stream_matmul_33_source_21_pat_size_1 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_count_2 <= _source_stream_matmul_33_source_21_pat_size_2 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_count_3 <= _source_stream_matmul_33_source_21_pat_size_3 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_size_buf_0 <= _source_stream_matmul_33_source_21_pat_size_0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_size_buf_1 <= _source_stream_matmul_33_source_21_pat_size_1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_size_buf_2 <= _source_stream_matmul_33_source_21_pat_size_2;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_size_buf_3 <= _source_stream_matmul_33_source_21_pat_size_3;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_stride_buf_0 <= _source_stream_matmul_33_source_21_pat_stride_0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_stride_buf_1 <= _source_stream_matmul_33_source_21_pat_stride_1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_stride_buf_2 <= _source_stream_matmul_33_source_21_pat_stride_2;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_stride_buf_3 <= _source_stream_matmul_33_source_21_pat_stride_3;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_source_busy && _stream_matmul_33_is_root) begin
        __variable_wdata_1158 <= _stream_matmul_33_source_21_source_ram_rdata;
      end 
      if((_stream_matmul_33_source_21_source_pat_fsm_3 == 1) && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_21_idle <= 0;
        _stream_matmul_33_source_21_source_ram_raddr <= _stream_matmul_33_source_21_source_pat_all_offset;
        _stream_matmul_33_source_21_source_ram_renable <= 1;
      end 
      if((_stream_matmul_33_source_21_source_pat_fsm_3 == 1) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_cur_offset_0 <= _source_stream_matmul_33_source_21_pat_cur_offset_0 + _source_stream_matmul_33_source_21_pat_stride_buf_0;
        _source_stream_matmul_33_source_21_pat_count_0 <= _source_stream_matmul_33_source_21_pat_count_0 - 1;
      end 
      if((_stream_matmul_33_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_33_source_21_pat_count_0 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_cur_offset_0 <= 0;
        _source_stream_matmul_33_source_21_pat_count_0 <= _source_stream_matmul_33_source_21_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_33_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_33_source_21_pat_count_0 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_cur_offset_1 <= _source_stream_matmul_33_source_21_pat_cur_offset_1 + _source_stream_matmul_33_source_21_pat_stride_buf_1;
        _source_stream_matmul_33_source_21_pat_count_1 <= _source_stream_matmul_33_source_21_pat_count_1 - 1;
      end 
      if((_stream_matmul_33_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_33_source_21_pat_count_0 == 0) && (_source_stream_matmul_33_source_21_pat_count_1 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_cur_offset_1 <= 0;
        _source_stream_matmul_33_source_21_pat_count_1 <= _source_stream_matmul_33_source_21_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_33_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_33_source_21_pat_count_0 == 0) && (_source_stream_matmul_33_source_21_pat_count_1 == 0)) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_cur_offset_2 <= _source_stream_matmul_33_source_21_pat_cur_offset_2 + _source_stream_matmul_33_source_21_pat_stride_buf_2;
        _source_stream_matmul_33_source_21_pat_count_2 <= _source_stream_matmul_33_source_21_pat_count_2 - 1;
      end 
      if((_stream_matmul_33_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_33_source_21_pat_count_0 == 0) && (_source_stream_matmul_33_source_21_pat_count_1 == 0)) && (_source_stream_matmul_33_source_21_pat_count_2 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_cur_offset_2 <= 0;
        _source_stream_matmul_33_source_21_pat_count_2 <= _source_stream_matmul_33_source_21_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_33_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_33_source_21_pat_count_0 == 0) && (_source_stream_matmul_33_source_21_pat_count_1 == 0) && (_source_stream_matmul_33_source_21_pat_count_2 == 0)) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_cur_offset_3 <= _source_stream_matmul_33_source_21_pat_cur_offset_3 + _source_stream_matmul_33_source_21_pat_stride_buf_3;
        _source_stream_matmul_33_source_21_pat_count_3 <= _source_stream_matmul_33_source_21_pat_count_3 - 1;
      end 
      if((_stream_matmul_33_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_33_source_21_pat_count_0 == 0) && (_source_stream_matmul_33_source_21_pat_count_1 == 0) && (_source_stream_matmul_33_source_21_pat_count_2 == 0)) && (_source_stream_matmul_33_source_21_pat_count_3 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_21_pat_cur_offset_3 <= 0;
        _source_stream_matmul_33_source_21_pat_count_3 <= _source_stream_matmul_33_source_21_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_33_source_21_source_pat_fsm_3 == 1) && _stream_matmul_33_source_stop && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_21_source_ram_renable <= 0;
        _stream_matmul_33_source_21_idle <= 1;
      end 
      if((_stream_matmul_33_source_21_source_pat_fsm_3 == 2) && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_21_source_ram_renable <= 0;
        _stream_matmul_33_source_21_idle <= 1;
      end 
      if(_set_flag_1699) begin
        _stream_matmul_33_source_22_source_mode <= 5'b10;
        _stream_matmul_33_source_22_source_offset <= matmul_33_filter_page_comp_offset_buf;
      end 
      if(_set_flag_1699) begin
        _source_stream_matmul_33_source_22_pat_size_0 <= cparam_matmul_33_stream_reduce_size;
        _source_stream_matmul_33_source_22_pat_stride_0 <= 1;
      end 
      if(_set_flag_1699) begin
        _source_stream_matmul_33_source_22_pat_size_1 <= matmul_33_next_stream_num_ops;
        _source_stream_matmul_33_source_22_pat_stride_1 <= cparam_matmul_33_stream_aligned_reduce_size;
      end 
      if(_set_flag_1699) begin
        _source_stream_matmul_33_source_22_pat_size_2 <= 1;
        _source_stream_matmul_33_source_22_pat_stride_2 <= 0;
      end 
      if(_set_flag_1699) begin
        _source_stream_matmul_33_source_22_pat_size_3 <= 1;
        _source_stream_matmul_33_source_22_pat_stride_3 <= 0;
      end 
      if(_set_flag_1699) begin
        _stream_matmul_33_source_22_source_sel <= 5;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_22_source_offset_buf <= _stream_matmul_33_source_22_source_offset;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_count_0 <= _source_stream_matmul_33_source_22_pat_size_0 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_count_1 <= _source_stream_matmul_33_source_22_pat_size_1 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_count_2 <= _source_stream_matmul_33_source_22_pat_size_2 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_count_3 <= _source_stream_matmul_33_source_22_pat_size_3 - 1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_size_buf_0 <= _source_stream_matmul_33_source_22_pat_size_0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_size_buf_1 <= _source_stream_matmul_33_source_22_pat_size_1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_size_buf_2 <= _source_stream_matmul_33_source_22_pat_size_2;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_size_buf_3 <= _source_stream_matmul_33_source_22_pat_size_3;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_stride_buf_0 <= _source_stream_matmul_33_source_22_pat_stride_0;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_stride_buf_1 <= _source_stream_matmul_33_source_22_pat_stride_1;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_stride_buf_2 <= _source_stream_matmul_33_source_22_pat_stride_2;
      end 
      if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_stride_buf_3 <= _source_stream_matmul_33_source_22_pat_stride_3;
      end 
      if(_stream_matmul_33_stream_oready && _stream_matmul_33_source_busy && _stream_matmul_33_is_root) begin
        __variable_wdata_1159 <= _stream_matmul_33_source_22_source_ram_rdata;
      end 
      if((_stream_matmul_33_source_22_source_pat_fsm_4 == 1) && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_22_idle <= 0;
        _stream_matmul_33_source_22_source_ram_raddr <= _stream_matmul_33_source_22_source_pat_all_offset;
        _stream_matmul_33_source_22_source_ram_renable <= 1;
      end 
      if((_stream_matmul_33_source_22_source_pat_fsm_4 == 1) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_cur_offset_0 <= _source_stream_matmul_33_source_22_pat_cur_offset_0 + _source_stream_matmul_33_source_22_pat_stride_buf_0;
        _source_stream_matmul_33_source_22_pat_count_0 <= _source_stream_matmul_33_source_22_pat_count_0 - 1;
      end 
      if((_stream_matmul_33_source_22_source_pat_fsm_4 == 1) && (_source_stream_matmul_33_source_22_pat_count_0 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_cur_offset_0 <= 0;
        _source_stream_matmul_33_source_22_pat_count_0 <= _source_stream_matmul_33_source_22_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_33_source_22_source_pat_fsm_4 == 1) && (_source_stream_matmul_33_source_22_pat_count_0 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_cur_offset_1 <= _source_stream_matmul_33_source_22_pat_cur_offset_1 + _source_stream_matmul_33_source_22_pat_stride_buf_1;
        _source_stream_matmul_33_source_22_pat_count_1 <= _source_stream_matmul_33_source_22_pat_count_1 - 1;
      end 
      if((_stream_matmul_33_source_22_source_pat_fsm_4 == 1) && (_source_stream_matmul_33_source_22_pat_count_0 == 0) && (_source_stream_matmul_33_source_22_pat_count_1 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_cur_offset_1 <= 0;
        _source_stream_matmul_33_source_22_pat_count_1 <= _source_stream_matmul_33_source_22_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_33_source_22_source_pat_fsm_4 == 1) && ((_source_stream_matmul_33_source_22_pat_count_0 == 0) && (_source_stream_matmul_33_source_22_pat_count_1 == 0)) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_cur_offset_2 <= _source_stream_matmul_33_source_22_pat_cur_offset_2 + _source_stream_matmul_33_source_22_pat_stride_buf_2;
        _source_stream_matmul_33_source_22_pat_count_2 <= _source_stream_matmul_33_source_22_pat_count_2 - 1;
      end 
      if((_stream_matmul_33_source_22_source_pat_fsm_4 == 1) && ((_source_stream_matmul_33_source_22_pat_count_0 == 0) && (_source_stream_matmul_33_source_22_pat_count_1 == 0)) && (_source_stream_matmul_33_source_22_pat_count_2 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_cur_offset_2 <= 0;
        _source_stream_matmul_33_source_22_pat_count_2 <= _source_stream_matmul_33_source_22_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_33_source_22_source_pat_fsm_4 == 1) && ((_source_stream_matmul_33_source_22_pat_count_0 == 0) && (_source_stream_matmul_33_source_22_pat_count_1 == 0) && (_source_stream_matmul_33_source_22_pat_count_2 == 0)) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_cur_offset_3 <= _source_stream_matmul_33_source_22_pat_cur_offset_3 + _source_stream_matmul_33_source_22_pat_stride_buf_3;
        _source_stream_matmul_33_source_22_pat_count_3 <= _source_stream_matmul_33_source_22_pat_count_3 - 1;
      end 
      if((_stream_matmul_33_source_22_source_pat_fsm_4 == 1) && ((_source_stream_matmul_33_source_22_pat_count_0 == 0) && (_source_stream_matmul_33_source_22_pat_count_1 == 0) && (_source_stream_matmul_33_source_22_pat_count_2 == 0)) && (_source_stream_matmul_33_source_22_pat_count_3 == 0) && _stream_matmul_33_stream_oready) begin
        _source_stream_matmul_33_source_22_pat_cur_offset_3 <= 0;
        _source_stream_matmul_33_source_22_pat_count_3 <= _source_stream_matmul_33_source_22_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_33_source_22_source_pat_fsm_4 == 1) && _stream_matmul_33_source_stop && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_22_source_ram_renable <= 0;
        _stream_matmul_33_source_22_idle <= 1;
      end 
      if((_stream_matmul_33_source_22_source_pat_fsm_4 == 2) && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_source_22_source_ram_renable <= 0;
        _stream_matmul_33_source_22_idle <= 1;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1703 <= _set_flag_1702;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1704 <= _tmp_1703;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1705 <= _tmp_1704;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1706 <= _tmp_1705;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1707 <= _tmp_1706;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1708 <= _tmp_1707;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1709 <= _tmp_1708;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1710 <= _tmp_1709;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1711 <= _tmp_1710;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1712 <= _tmp_1711;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1713 <= _tmp_1712;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1714 <= _tmp_1713;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1715 <= _tmp_1714;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1716 <= _tmp_1715;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1717 <= _tmp_1716;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1718 <= _tmp_1717;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1719 <= _tmp_1718;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1720 <= _tmp_1719;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1721 <= _tmp_1720;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1722 <= _tmp_1721;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1723 <= _tmp_1722;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1724 <= _tmp_1723;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1725 <= _tmp_1724;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1726 <= _tmp_1725;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1727 <= _tmp_1726;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1728 <= _tmp_1727;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1729 <= _tmp_1728;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1730 <= _tmp_1729;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1731 <= _tmp_1730;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1732 <= _tmp_1731;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1733 <= _tmp_1732;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1734 <= _tmp_1733;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1737 <= _tmp_1736;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1738 <= _tmp_1737;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1739 <= _tmp_1738;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1740 <= _tmp_1739;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1741 <= _tmp_1740;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1742 <= _tmp_1741;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1743 <= _tmp_1742;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1744 <= _tmp_1743;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1745 <= _tmp_1744;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1746 <= _tmp_1745;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1747 <= _tmp_1746;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1748 <= _tmp_1747;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1749 <= _tmp_1748;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1750 <= _tmp_1749;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1751 <= _tmp_1750;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1752 <= _tmp_1751;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1753 <= _tmp_1752;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1754 <= _tmp_1753;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1755 <= _tmp_1754;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1756 <= _tmp_1755;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1757 <= _tmp_1756;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1758 <= _tmp_1757;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1759 <= _tmp_1758;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1760 <= _tmp_1759;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1761 <= _tmp_1760;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1762 <= _tmp_1761;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1763 <= _tmp_1762;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1764 <= _tmp_1763;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1765 <= _tmp_1764;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1766 <= _tmp_1765;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1767 <= _tmp_1766;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1768 <= _tmp_1767;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1769 <= matmul_33_next_stream_num_ops;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1770 <= _tmp_1769;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1771 <= _tmp_1770;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1772 <= _tmp_1771;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1773 <= _tmp_1772;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1774 <= _tmp_1773;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1775 <= _tmp_1774;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1776 <= _tmp_1775;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1777 <= _tmp_1776;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1778 <= _tmp_1777;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1779 <= _tmp_1778;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1780 <= _tmp_1779;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1781 <= _tmp_1780;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1782 <= _tmp_1781;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1783 <= _tmp_1782;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1784 <= _tmp_1783;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1785 <= _tmp_1784;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1786 <= _tmp_1785;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1787 <= _tmp_1786;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1788 <= _tmp_1787;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1789 <= _tmp_1788;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1790 <= _tmp_1789;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1791 <= _tmp_1790;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1792 <= _tmp_1791;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1793 <= _tmp_1792;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1794 <= _tmp_1793;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1795 <= _tmp_1794;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1796 <= _tmp_1795;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1797 <= _tmp_1796;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1798 <= _tmp_1797;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1799 <= _tmp_1798;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1800 <= _tmp_1799;
      end 
      if(_tmp_1734) begin
        _stream_matmul_33_sink_33_sink_mode <= 5'b1;
        _stream_matmul_33_sink_33_sink_offset <= _tmp_1768;
        _stream_matmul_33_sink_33_sink_size <= _tmp_1800;
        _stream_matmul_33_sink_33_sink_stride <= 1;
      end 
      if(_tmp_1734) begin
        _stream_matmul_33_sink_33_sink_sel <= 6;
      end 
      if(_stream_matmul_33_sink_start && _stream_matmul_33_sink_33_sink_mode & 5'b1 && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_sink_33_sink_offset_buf <= _stream_matmul_33_sink_33_sink_offset;
        _stream_matmul_33_sink_33_sink_size_buf <= _stream_matmul_33_sink_33_sink_size;
        _stream_matmul_33_sink_33_sink_stride_buf <= _stream_matmul_33_sink_33_sink_stride;
      end 
      if((_stream_matmul_33_sink_33_sink_fsm_5 == 1) && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_sink_33_sink_waddr <= _stream_matmul_33_sink_33_sink_offset_buf - _stream_matmul_33_sink_33_sink_stride_buf;
        _stream_matmul_33_sink_33_sink_count <= _stream_matmul_33_sink_33_sink_size_buf;
      end 
      if((_stream_matmul_33_sink_33_sink_fsm_5 == 2) && stream_matmul_33_sink_34_data && _stream_matmul_33_stream_oready) begin
        _stream_matmul_33_sink_33_sink_waddr <= _stream_matmul_33_sink_33_sink_waddr + _stream_matmul_33_sink_33_sink_stride_buf;
        _stream_matmul_33_sink_33_sink_wdata <= stream_matmul_33_sink_33_data;
        _stream_matmul_33_sink_33_sink_wenable <= 1;
        _stream_matmul_33_sink_33_sink_count <= _stream_matmul_33_sink_33_sink_count - 1;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1894 <= _stream_matmul_33_source_start;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1895 <= _tmp_1894;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1896 <= _tmp_1895;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1897 <= _stream_matmul_33_source_start;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1898 <= _tmp_1897;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1899 <= _tmp_1898;
      end 
      if(_stream_matmul_33_stream_oready && _tmp_1899) begin
        __variable_wdata_1057 <= 1;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1900 <= _stream_matmul_33_source_start;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1901 <= _tmp_1900;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1902 <= _tmp_1901;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1903 <= _tmp_1902;
      end 
      if(_stream_matmul_33_stream_oready && _tmp_1903) begin
        __variable_wdata_1057 <= 0;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1906 <= _tmp_1905;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1909 <= _tmp_1908;
      end 
      if(_stream_matmul_33_stream_oready && _tmp_1909) begin
        __variable_wdata_1057 <= 1;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1910 <= _stream_matmul_33_source_start;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1911 <= _tmp_1910;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1912 <= _tmp_1911;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1913 <= _tmp_1912;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1914 <= _tmp_1913;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1915 <= _tmp_1914;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1916 <= _tmp_1915;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1917 <= _tmp_1916;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1918 <= _tmp_1917;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1919 <= _tmp_1918;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1920 <= _tmp_1919;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1921 <= _tmp_1920;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1922 <= _tmp_1921;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1923 <= _tmp_1922;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1924 <= _tmp_1923;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1925 <= _tmp_1924;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1926 <= _tmp_1925;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1927 <= _tmp_1926;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1928 <= _tmp_1927;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1929 <= _tmp_1928;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1930 <= _tmp_1929;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1931 <= _tmp_1930;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1932 <= _tmp_1931;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1933 <= _tmp_1932;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1934 <= _tmp_1933;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1935 <= _tmp_1934;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1936 <= _tmp_1935;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1937 <= _tmp_1936;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1938 <= _tmp_1937;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1939 <= _tmp_1938;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1940 <= _tmp_1939;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1941 <= _tmp_1940;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1942 <= _stream_matmul_33_source_stop;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1943 <= _tmp_1942;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1944 <= _tmp_1943;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1945 <= _tmp_1944;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1946 <= _tmp_1945;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1947 <= _tmp_1946;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1948 <= _tmp_1947;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1949 <= _tmp_1948;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1950 <= _tmp_1949;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1951 <= _tmp_1950;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1952 <= _tmp_1951;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1953 <= _tmp_1952;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1954 <= _tmp_1953;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1955 <= _tmp_1954;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1956 <= _tmp_1955;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1957 <= _tmp_1956;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1958 <= _tmp_1957;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1959 <= _tmp_1958;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1960 <= _tmp_1959;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1961 <= _tmp_1960;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1962 <= _tmp_1961;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1963 <= _tmp_1962;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1964 <= _tmp_1963;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1965 <= _tmp_1964;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1966 <= _tmp_1965;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1967 <= _tmp_1966;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1968 <= _tmp_1967;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1969 <= _tmp_1968;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1970 <= _tmp_1969;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1971 <= _tmp_1970;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1972 <= _tmp_1971;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1973 <= _tmp_1972;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1974 <= _stream_matmul_33_source_busy;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1975 <= _tmp_1974;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1976 <= _tmp_1975;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1977 <= _tmp_1976;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1978 <= _tmp_1977;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1979 <= _tmp_1978;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1980 <= _tmp_1979;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1981 <= _tmp_1980;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1982 <= _tmp_1981;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1983 <= _tmp_1982;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1984 <= _tmp_1983;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1985 <= _tmp_1984;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1986 <= _tmp_1985;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1987 <= _tmp_1986;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1988 <= _tmp_1987;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1989 <= _tmp_1988;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1990 <= _tmp_1989;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1991 <= _tmp_1990;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1992 <= _tmp_1991;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1993 <= _tmp_1992;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1994 <= _tmp_1993;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1995 <= _tmp_1994;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1996 <= _tmp_1995;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1997 <= _tmp_1996;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1998 <= _tmp_1997;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_1999 <= _tmp_1998;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_2000 <= _tmp_1999;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_2001 <= _tmp_2000;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_2002 <= _tmp_2001;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_2003 <= _tmp_2002;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_2004 <= _tmp_2003;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_2005 <= _tmp_2004;
      end 
      if(_stream_matmul_33_stream_oready) begin
        _tmp_2006 <= _stream_matmul_33_sink_busy;
      end 
      if(!_stream_matmul_33_sink_busy && _tmp_2006) begin
        _stream_matmul_33_busy_reg <= 0;
      end 
      if(_stream_matmul_33_source_busy) begin
        _stream_matmul_33_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_matmul_33_fsm_1 = 1;
  localparam _stream_matmul_33_fsm_2 = 2;
  localparam _stream_matmul_33_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_33_fsm <= _stream_matmul_33_fsm_init;
      _stream_matmul_33_source_start <= 0;
      _stream_matmul_33_source_busy <= 0;
      _stream_matmul_33_stream_ivalid <= 0;
    end else begin
      if(_stream_matmul_33_stream_oready && _tmp_1896) begin
        _stream_matmul_33_stream_ivalid <= 1;
      end 
      if(_stream_matmul_33_stream_oready && _tmp_1906) begin
        _stream_matmul_33_stream_ivalid <= 0;
      end 
      case(_stream_matmul_33_fsm)
        _stream_matmul_33_fsm_init: begin
          if(_stream_matmul_33_run_flag) begin
            _stream_matmul_33_source_start <= 1;
          end 
          if(_stream_matmul_33_run_flag) begin
            _stream_matmul_33_fsm <= _stream_matmul_33_fsm_1;
          end 
        end
        _stream_matmul_33_fsm_1: begin
          if(_stream_matmul_33_source_start && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_start <= 0;
            _stream_matmul_33_source_busy <= 1;
          end 
          if(_stream_matmul_33_source_start && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_fsm <= _stream_matmul_33_fsm_2;
          end 
        end
        _stream_matmul_33_fsm_2: begin
          if(_stream_matmul_33_stream_oready) begin
            _stream_matmul_33_fsm <= _stream_matmul_33_fsm_3;
          end 
        end
        _stream_matmul_33_fsm_3: begin
          if(_stream_matmul_33_stream_oready && (_stream_matmul_33_source_11_idle && _stream_matmul_33_source_13_idle && _stream_matmul_33_source_15_idle && _stream_matmul_33_source_20_idle && _stream_matmul_33_source_21_idle && _stream_matmul_33_source_22_idle && _stream_matmul_33_source_7_idle && _stream_matmul_33_source_9_idle && (_stream_matmul_33_fsm == 3))) begin
            _stream_matmul_33_source_busy <= 0;
          end 
          if(_stream_matmul_33_stream_oready && (_stream_matmul_33_source_11_idle && _stream_matmul_33_source_13_idle && _stream_matmul_33_source_15_idle && _stream_matmul_33_source_20_idle && _stream_matmul_33_source_21_idle && _stream_matmul_33_source_22_idle && _stream_matmul_33_source_7_idle && _stream_matmul_33_source_9_idle && (_stream_matmul_33_fsm == 3)) && _stream_matmul_33_run_flag) begin
            _stream_matmul_33_source_start <= 1;
          end 
          if(_stream_matmul_33_stream_oready && (_stream_matmul_33_source_11_idle && _stream_matmul_33_source_13_idle && _stream_matmul_33_source_15_idle && _stream_matmul_33_source_20_idle && _stream_matmul_33_source_21_idle && _stream_matmul_33_source_22_idle && _stream_matmul_33_source_7_idle && _stream_matmul_33_source_9_idle && (_stream_matmul_33_fsm == 3))) begin
            _stream_matmul_33_fsm <= _stream_matmul_33_fsm_init;
          end 
          if(_stream_matmul_33_stream_oready && (_stream_matmul_33_source_11_idle && _stream_matmul_33_source_13_idle && _stream_matmul_33_source_15_idle && _stream_matmul_33_source_20_idle && _stream_matmul_33_source_21_idle && _stream_matmul_33_source_22_idle && _stream_matmul_33_source_7_idle && _stream_matmul_33_source_9_idle && (_stream_matmul_33_fsm == 3)) && _stream_matmul_33_run_flag) begin
            _stream_matmul_33_fsm <= _stream_matmul_33_fsm_1;
          end 
        end
      endcase
    end
  end

  localparam main_fsm_1 = 1;
  localparam main_fsm_2 = 2;
  localparam main_fsm_3 = 3;
  localparam main_fsm_4 = 4;
  localparam main_fsm_5 = 5;
  localparam main_fsm_6 = 6;
  localparam main_fsm_7 = 7;
  localparam main_fsm_8 = 8;
  localparam main_fsm_9 = 9;
  localparam main_fsm_10 = 10;
  localparam main_fsm_11 = 11;
  localparam main_fsm_12 = 12;
  localparam main_fsm_13 = 13;
  localparam main_fsm_14 = 14;
  localparam main_fsm_15 = 15;
  localparam main_fsm_16 = 16;
  localparam main_fsm_17 = 17;
  localparam main_fsm_18 = 18;
  localparam main_fsm_19 = 19;
  localparam main_fsm_20 = 20;
  localparam main_fsm_21 = 21;
  localparam main_fsm_22 = 22;
  localparam main_fsm_23 = 23;
  localparam main_fsm_24 = 24;
  localparam main_fsm_25 = 25;
  localparam main_fsm_26 = 26;
  localparam main_fsm_27 = 27;
  localparam main_fsm_28 = 28;
  localparam main_fsm_29 = 29;
  localparam main_fsm_30 = 30;
  localparam main_fsm_31 = 31;
  localparam main_fsm_32 = 32;
  localparam main_fsm_33 = 33;
  localparam main_fsm_34 = 34;
  localparam main_fsm_35 = 35;
  localparam main_fsm_36 = 36;
  localparam main_fsm_37 = 37;
  localparam main_fsm_38 = 38;
  localparam main_fsm_39 = 39;
  localparam main_fsm_40 = 40;
  localparam main_fsm_41 = 41;
  localparam main_fsm_42 = 42;
  localparam main_fsm_43 = 43;
  localparam main_fsm_44 = 44;
  localparam main_fsm_45 = 45;
  localparam main_fsm_46 = 46;
  localparam main_fsm_47 = 47;
  localparam main_fsm_48 = 48;
  localparam main_fsm_49 = 49;
  localparam main_fsm_50 = 50;
  localparam main_fsm_51 = 51;
  localparam main_fsm_52 = 52;
  localparam main_fsm_53 = 53;
  localparam main_fsm_54 = 54;
  localparam main_fsm_55 = 55;
  localparam main_fsm_56 = 56;
  localparam main_fsm_57 = 57;
  localparam main_fsm_58 = 58;
  localparam main_fsm_59 = 59;
  localparam main_fsm_60 = 60;
  localparam main_fsm_61 = 61;
  localparam main_fsm_62 = 62;
  localparam main_fsm_63 = 63;
  localparam main_fsm_64 = 64;
  localparam main_fsm_65 = 65;
  localparam main_fsm_66 = 66;
  localparam main_fsm_67 = 67;
  localparam main_fsm_68 = 68;
  localparam main_fsm_69 = 69;
  localparam main_fsm_70 = 70;
  localparam main_fsm_71 = 71;
  localparam main_fsm_72 = 72;
  localparam main_fsm_73 = 73;
  localparam main_fsm_74 = 74;
  localparam main_fsm_75 = 75;
  localparam main_fsm_76 = 76;
  localparam main_fsm_77 = 77;
  localparam main_fsm_78 = 78;
  localparam main_fsm_79 = 79;
  localparam main_fsm_80 = 80;
  localparam main_fsm_81 = 81;
  localparam main_fsm_82 = 82;
  localparam main_fsm_83 = 83;
  localparam main_fsm_84 = 84;
  localparam main_fsm_85 = 85;
  localparam main_fsm_86 = 86;
  localparam main_fsm_87 = 87;
  localparam main_fsm_88 = 88;
  localparam main_fsm_89 = 89;
  localparam main_fsm_90 = 90;
  localparam main_fsm_91 = 91;

  always @(posedge CLK) begin
    if(RST) begin
      main_fsm <= main_fsm_init;
      conv2d_4_objaddr <= 0;
      conv2d_4_arg_objaddr_0 <= 0;
      conv2d_4_arg_objaddr_1 <= 0;
      conv2d_4_arg_objaddr_2 <= 0;
      conv2d_4_arg_objaddr_3 <= 0;
      conv2d_4_control_param_index <= 0;
      max_pool_serial_6_objaddr <= 0;
      max_pool_serial_6_arg_objaddr_0 <= 0;
      max_pool_serial_6_control_param_index <= 0;
      matmul_23_objaddr <= 0;
      matmul_23_arg_objaddr_0 <= 0;
      matmul_23_arg_objaddr_1 <= 0;
      matmul_23_arg_objaddr_2 <= 0;
      matmul_23_arg_objaddr_3 <= 0;
      matmul_23_control_param_index <= 0;
      matmul_33_objaddr <= 0;
      matmul_33_arg_objaddr_0 <= 0;
      matmul_33_arg_objaddr_1 <= 0;
      matmul_33_arg_objaddr_2 <= 0;
      matmul_33_arg_objaddr_3 <= 0;
    end else begin
      case(main_fsm)
        main_fsm_init: begin
          if(_saxi_register_4 != 0) begin
            main_fsm <= main_fsm_1;
          end 
        end
        main_fsm_1: begin
          main_fsm <= main_fsm_2;
        end
        main_fsm_2: begin
          main_fsm <= main_fsm_3;
        end
        main_fsm_3: begin
          main_fsm <= main_fsm_4;
        end
        main_fsm_4: begin
          main_fsm <= main_fsm_5;
        end
        main_fsm_5: begin
          conv2d_4_objaddr <= _saxi_register_33;
          main_fsm <= main_fsm_6;
        end
        main_fsm_6: begin
          conv2d_4_arg_objaddr_0 <= _saxi_register_35;
          main_fsm <= main_fsm_7;
        end
        main_fsm_7: begin
          conv2d_4_arg_objaddr_1 <= _saxi_register_36;
          main_fsm <= main_fsm_8;
        end
        main_fsm_8: begin
          conv2d_4_arg_objaddr_2 <= _saxi_register_36 + 4608;
          main_fsm <= main_fsm_9;
        end
        main_fsm_9: begin
          conv2d_4_arg_objaddr_3 <= _saxi_register_36 + 4736;
          main_fsm <= main_fsm_10;
        end
        main_fsm_10: begin
          conv2d_4_control_param_index <= 0;
          main_fsm <= main_fsm_11;
        end
        main_fsm_11: begin
          main_fsm <= main_fsm_12;
        end
        main_fsm_12: begin
          main_fsm <= main_fsm_13;
        end
        main_fsm_13: begin
          if(control_conv2d_4 == 34) begin
            main_fsm <= main_fsm_14;
          end 
        end
        main_fsm_14: begin
          main_fsm <= main_fsm_15;
        end
        main_fsm_15: begin
          max_pool_serial_6_objaddr <= _saxi_register_33 + 131072;
          main_fsm <= main_fsm_16;
        end
        main_fsm_16: begin
          max_pool_serial_6_arg_objaddr_0 <= _saxi_register_33;
          main_fsm <= main_fsm_17;
        end
        main_fsm_17: begin
          max_pool_serial_6_control_param_index <= 0;
          main_fsm <= main_fsm_18;
        end
        main_fsm_18: begin
          main_fsm <= main_fsm_19;
        end
        main_fsm_19: begin
          main_fsm <= main_fsm_20;
        end
        main_fsm_20: begin
          if(control_max_pool_serial_6 == 19) begin
            main_fsm <= main_fsm_21;
          end 
        end
        main_fsm_21: begin
          main_fsm <= main_fsm_22;
        end
        main_fsm_22: begin
          conv2d_4_objaddr <= _saxi_register_33 + 163840;
          main_fsm <= main_fsm_23;
        end
        main_fsm_23: begin
          conv2d_4_arg_objaddr_0 <= _saxi_register_33 + 131072;
          main_fsm <= main_fsm_24;
        end
        main_fsm_24: begin
          conv2d_4_arg_objaddr_1 <= _saxi_register_36 + 4864;
          main_fsm <= main_fsm_25;
        end
        main_fsm_25: begin
          conv2d_4_arg_objaddr_2 <= _saxi_register_36 + 152320;
          main_fsm <= main_fsm_26;
        end
        main_fsm_26: begin
          conv2d_4_arg_objaddr_3 <= _saxi_register_36 + 152576;
          main_fsm <= main_fsm_27;
        end
        main_fsm_27: begin
          conv2d_4_control_param_index <= 1;
          main_fsm <= main_fsm_28;
        end
        main_fsm_28: begin
          main_fsm <= main_fsm_29;
        end
        main_fsm_29: begin
          main_fsm <= main_fsm_30;
        end
        main_fsm_30: begin
          if(control_conv2d_4 == 34) begin
            main_fsm <= main_fsm_31;
          end 
        end
        main_fsm_31: begin
          main_fsm <= main_fsm_32;
        end
        main_fsm_32: begin
          max_pool_serial_6_objaddr <= _saxi_register_33 + 229376;
          main_fsm <= main_fsm_33;
        end
        main_fsm_33: begin
          max_pool_serial_6_arg_objaddr_0 <= _saxi_register_33 + 163840;
          main_fsm <= main_fsm_34;
        end
        main_fsm_34: begin
          max_pool_serial_6_control_param_index <= 1;
          main_fsm <= main_fsm_35;
        end
        main_fsm_35: begin
          main_fsm <= main_fsm_36;
        end
        main_fsm_36: begin
          main_fsm <= main_fsm_37;
        end
        main_fsm_37: begin
          if(control_max_pool_serial_6 == 19) begin
            main_fsm <= main_fsm_38;
          end 
        end
        main_fsm_38: begin
          main_fsm <= main_fsm_39;
        end
        main_fsm_39: begin
          conv2d_4_objaddr <= _saxi_register_33 + 245760;
          main_fsm <= main_fsm_40;
        end
        main_fsm_40: begin
          conv2d_4_arg_objaddr_0 <= _saxi_register_33 + 229376;
          main_fsm <= main_fsm_41;
        end
        main_fsm_41: begin
          conv2d_4_arg_objaddr_1 <= _saxi_register_36 + 152832;
          main_fsm <= main_fsm_42;
        end
        main_fsm_42: begin
          conv2d_4_arg_objaddr_2 <= _saxi_register_36 + 742656;
          main_fsm <= main_fsm_43;
        end
        main_fsm_43: begin
          conv2d_4_arg_objaddr_3 <= _saxi_register_36 + 743168;
          main_fsm <= main_fsm_44;
        end
        main_fsm_44: begin
          conv2d_4_control_param_index <= 2;
          main_fsm <= main_fsm_45;
        end
        main_fsm_45: begin
          main_fsm <= main_fsm_46;
        end
        main_fsm_46: begin
          main_fsm <= main_fsm_47;
        end
        main_fsm_47: begin
          if(control_conv2d_4 == 34) begin
            main_fsm <= main_fsm_48;
          end 
        end
        main_fsm_48: begin
          main_fsm <= main_fsm_49;
        end
        main_fsm_49: begin
          max_pool_serial_6_objaddr <= _saxi_register_33 + 278528;
          main_fsm <= main_fsm_50;
        end
        main_fsm_50: begin
          max_pool_serial_6_arg_objaddr_0 <= _saxi_register_33 + 245760;
          main_fsm <= main_fsm_51;
        end
        main_fsm_51: begin
          max_pool_serial_6_control_param_index <= 2;
          main_fsm <= main_fsm_52;
        end
        main_fsm_52: begin
          main_fsm <= main_fsm_53;
        end
        main_fsm_53: begin
          main_fsm <= main_fsm_54;
        end
        main_fsm_54: begin
          if(control_max_pool_serial_6 == 19) begin
            main_fsm <= main_fsm_55;
          end 
        end
        main_fsm_55: begin
          main_fsm <= main_fsm_56;
        end
        main_fsm_56: begin
          main_fsm <= main_fsm_57;
        end
        main_fsm_57: begin
          main_fsm <= main_fsm_58;
        end
        main_fsm_58: begin
          matmul_23_objaddr <= _saxi_register_33 + 286720;
          main_fsm <= main_fsm_59;
        end
        main_fsm_59: begin
          matmul_23_arg_objaddr_0 <= _saxi_register_33 + 278528;
          main_fsm <= main_fsm_60;
        end
        main_fsm_60: begin
          matmul_23_arg_objaddr_1 <= _saxi_register_36 + 743680;
          main_fsm <= main_fsm_61;
        end
        main_fsm_61: begin
          matmul_23_arg_objaddr_2 <= _saxi_register_36 + 9132288;
          main_fsm <= main_fsm_62;
        end
        main_fsm_62: begin
          matmul_23_arg_objaddr_3 <= _saxi_register_36 + 9134336;
          main_fsm <= main_fsm_63;
        end
        main_fsm_63: begin
          matmul_23_control_param_index <= 0;
          main_fsm <= main_fsm_64;
        end
        main_fsm_64: begin
          main_fsm <= main_fsm_65;
        end
        main_fsm_65: begin
          main_fsm <= main_fsm_66;
        end
        main_fsm_66: begin
          if(control_matmul_23 == 28) begin
            main_fsm <= main_fsm_67;
          end 
        end
        main_fsm_67: begin
          main_fsm <= main_fsm_68;
        end
        main_fsm_68: begin
          matmul_23_objaddr <= _saxi_register_33 + 288768;
          main_fsm <= main_fsm_69;
        end
        main_fsm_69: begin
          matmul_23_arg_objaddr_0 <= _saxi_register_33 + 286720;
          main_fsm <= main_fsm_70;
        end
        main_fsm_70: begin
          matmul_23_arg_objaddr_1 <= _saxi_register_36 + 9136384;
          main_fsm <= main_fsm_71;
        end
        main_fsm_71: begin
          matmul_23_arg_objaddr_2 <= _saxi_register_36 + 10184960;
          main_fsm <= main_fsm_72;
        end
        main_fsm_72: begin
          matmul_23_arg_objaddr_3 <= _saxi_register_36 + 10185984;
          main_fsm <= main_fsm_73;
        end
        main_fsm_73: begin
          matmul_23_control_param_index <= 1;
          main_fsm <= main_fsm_74;
        end
        main_fsm_74: begin
          main_fsm <= main_fsm_75;
        end
        main_fsm_75: begin
          main_fsm <= main_fsm_76;
        end
        main_fsm_76: begin
          if(control_matmul_23 == 28) begin
            main_fsm <= main_fsm_77;
          end 
        end
        main_fsm_77: begin
          main_fsm <= main_fsm_78;
        end
        main_fsm_78: begin
          matmul_33_objaddr <= _saxi_register_34;
          main_fsm <= main_fsm_79;
        end
        main_fsm_79: begin
          matmul_33_arg_objaddr_0 <= _saxi_register_33 + 288768;
          main_fsm <= main_fsm_80;
        end
        main_fsm_80: begin
          matmul_33_arg_objaddr_1 <= _saxi_register_36 + 10187008;
          main_fsm <= main_fsm_81;
        end
        main_fsm_81: begin
          matmul_33_arg_objaddr_2 <= _saxi_register_36 + 10197248;
          main_fsm <= main_fsm_82;
        end
        main_fsm_82: begin
          matmul_33_arg_objaddr_3 <= _saxi_register_36 + 10197312;
          main_fsm <= main_fsm_83;
        end
        main_fsm_83: begin
          main_fsm <= main_fsm_84;
        end
        main_fsm_84: begin
          main_fsm <= main_fsm_85;
        end
        main_fsm_85: begin
          if(control_matmul_33 == 28) begin
            main_fsm <= main_fsm_86;
          end 
        end
        main_fsm_86: begin
          main_fsm <= main_fsm_87;
        end
        main_fsm_87: begin
          main_fsm <= main_fsm_88;
        end
        main_fsm_88: begin
          main_fsm <= main_fsm_89;
        end
        main_fsm_89: begin
          main_fsm <= main_fsm_90;
        end
        main_fsm_90: begin
          main_fsm <= main_fsm_91;
        end
        main_fsm_91: begin
          main_fsm <= main_fsm_init;
        end
      endcase
    end
  end

  localparam control_conv2d_4_1 = 1;
  localparam control_conv2d_4_2 = 2;
  localparam control_conv2d_4_3 = 3;
  localparam control_conv2d_4_4 = 4;
  localparam control_conv2d_4_5 = 5;
  localparam control_conv2d_4_6 = 6;
  localparam control_conv2d_4_7 = 7;
  localparam control_conv2d_4_8 = 8;
  localparam control_conv2d_4_9 = 9;
  localparam control_conv2d_4_10 = 10;
  localparam control_conv2d_4_11 = 11;
  localparam control_conv2d_4_12 = 12;
  localparam control_conv2d_4_13 = 13;
  localparam control_conv2d_4_14 = 14;
  localparam control_conv2d_4_15 = 15;
  localparam control_conv2d_4_16 = 16;
  localparam control_conv2d_4_17 = 17;
  localparam control_conv2d_4_18 = 18;
  localparam control_conv2d_4_19 = 19;
  localparam control_conv2d_4_20 = 20;
  localparam control_conv2d_4_21 = 21;
  localparam control_conv2d_4_22 = 22;
  localparam control_conv2d_4_23 = 23;
  localparam control_conv2d_4_24 = 24;
  localparam control_conv2d_4_25 = 25;
  localparam control_conv2d_4_26 = 26;
  localparam control_conv2d_4_27 = 27;
  localparam control_conv2d_4_28 = 28;
  localparam control_conv2d_4_29 = 29;
  localparam control_conv2d_4_30 = 30;
  localparam control_conv2d_4_31 = 31;
  localparam control_conv2d_4_32 = 32;
  localparam control_conv2d_4_33 = 33;
  localparam control_conv2d_4_34 = 34;

  always @(posedge CLK) begin
    if(RST) begin
      control_conv2d_4 <= control_conv2d_4_init;
      _control_conv2d_4_called <= 0;
      conv2d_4_filter_base_offset <= 0;
      conv2d_4_filter_page_comp_offset <= 0;
      conv2d_4_filter_page_dma_offset <= 0;
      conv2d_4_act_base_offset_row <= 0;
      conv2d_4_act_base_offset_bat <= 0;
      conv2d_4_dma_flag_0 <= 0;
      conv2d_4_dma_flag_1 <= 0;
      conv2d_4_dma_flag_2 <= 0;
      conv2d_4_act_page_comp_offset_0 <= 0;
      conv2d_4_act_page_comp_offset_1 <= 0;
      conv2d_4_act_page_comp_offset_2 <= 0;
      conv2d_4_act_page_dma_offset_0 <= 0;
      conv2d_4_act_page_dma_offset_1 <= 0;
      conv2d_4_act_page_dma_offset_2 <= 0;
      conv2d_4_out_base_offset_val <= 0;
      conv2d_4_out_base_offset_col <= 0;
      conv2d_4_out_base_offset_row <= 0;
      conv2d_4_out_base_offset_bat <= 0;
      conv2d_4_out_base_offset_och <= 0;
      conv2d_4_out_page <= 0;
      conv2d_4_out_page_comp_offset <= 0;
      conv2d_4_out_page_dma_offset <= 0;
      conv2d_4_out_laddr_offset <= 0;
      conv2d_4_sync_out_count <= 0;
      conv2d_4_write_count <= 0;
      conv2d_4_next_out_write_size <= 0;
      conv2d_4_row_count <= 0;
      conv2d_4_bat_count <= 0;
      conv2d_4_och_count <= 0;
      conv2d_4_row_select <= 0;
      conv2d_4_prev_row_count <= 0;
      conv2d_4_prev_bat_count <= 0;
      conv2d_4_prev_och_count <= 0;
      conv2d_4_prev_row_select <= 0;
      conv2d_4_out_col_count <= 0;
      conv2d_4_out_row_count <= 0;
      conv2d_4_out_ram_select <= 0;
      conv2d_4_skip_read_filter <= 0;
      conv2d_4_skip_read_act <= 0;
      conv2d_4_skip_comp <= 0;
      conv2d_4_skip_write_out <= 1;
    end else begin
      case(control_conv2d_4)
        control_conv2d_4_init: begin
          if(main_fsm == 11) begin
            _control_conv2d_4_called <= 1;
          end 
          if(main_fsm == 28) begin
            _control_conv2d_4_called <= 1;
          end 
          if(main_fsm == 45) begin
            _control_conv2d_4_called <= 1;
          end 
          if(main_fsm == 11) begin
            control_conv2d_4 <= control_conv2d_4_1;
          end 
          if(main_fsm == 28) begin
            control_conv2d_4 <= control_conv2d_4_1;
          end 
          if(main_fsm == 45) begin
            control_conv2d_4 <= control_conv2d_4_1;
          end 
        end
        control_conv2d_4_1: begin
          control_conv2d_4 <= control_conv2d_4_2;
        end
        control_conv2d_4_2: begin
          conv2d_4_filter_base_offset <= 0;
          conv2d_4_filter_page_comp_offset <= 0;
          conv2d_4_filter_page_dma_offset <= 0;
          conv2d_4_act_base_offset_row <= 0;
          conv2d_4_act_base_offset_bat <= 0;
          conv2d_4_dma_flag_0 <= 1;
          conv2d_4_dma_flag_1 <= 1;
          conv2d_4_dma_flag_2 <= 1;
          conv2d_4_act_page_comp_offset_0 <= 0;
          conv2d_4_act_page_comp_offset_1 <= 0;
          conv2d_4_act_page_comp_offset_2 <= 0;
          conv2d_4_act_page_dma_offset_0 <= 0;
          conv2d_4_act_page_dma_offset_1 <= 0;
          conv2d_4_act_page_dma_offset_2 <= 0;
          conv2d_4_out_base_offset_val <= 0;
          conv2d_4_out_base_offset_col <= 0;
          conv2d_4_out_base_offset_row <= 0;
          conv2d_4_out_base_offset_bat <= 0;
          conv2d_4_out_base_offset_och <= 0;
          conv2d_4_out_page <= 0;
          conv2d_4_out_page_comp_offset <= 0;
          conv2d_4_out_page_dma_offset <= 0;
          conv2d_4_out_laddr_offset <= 0;
          conv2d_4_sync_out_count <= 0;
          conv2d_4_write_count <= 0;
          conv2d_4_next_out_write_size <= (cparam_conv2d_4_max_och_count == 0)? cparam_conv2d_4_out_write_size_res : cparam_conv2d_4_out_write_size;
          conv2d_4_row_count <= 0;
          conv2d_4_bat_count <= 0;
          conv2d_4_och_count <= 0;
          conv2d_4_row_select <= 0;
          conv2d_4_prev_row_count <= 0;
          conv2d_4_prev_bat_count <= 0;
          conv2d_4_prev_och_count <= 0;
          conv2d_4_prev_row_select <= 0;
          conv2d_4_out_col_count <= 0;
          conv2d_4_out_row_count <= 0;
          conv2d_4_out_ram_select <= 0;
          conv2d_4_skip_read_filter <= 0;
          conv2d_4_skip_read_act <= 0;
          conv2d_4_skip_comp <= 0;
          conv2d_4_skip_write_out <= 1;
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_3;
          end 
        end
        control_conv2d_4_3: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_4;
          end 
        end
        control_conv2d_4_4: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_5;
          end 
        end
        control_conv2d_4_5: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_6;
          end 
        end
        control_conv2d_4_6: begin
          if(cparam_conv2d_4_data_stationary == 0) begin
            control_conv2d_4 <= control_conv2d_4_7;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            control_conv2d_4 <= control_conv2d_4_12;
          end 
        end
        control_conv2d_4_7: begin
          control_conv2d_4 <= control_conv2d_4_8;
          if(conv2d_4_skip_read_filter) begin
            control_conv2d_4 <= control_conv2d_4_11;
          end 
        end
        control_conv2d_4_8: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_9;
          end 
        end
        control_conv2d_4_9: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_10;
          end 
        end
        control_conv2d_4_10: begin
          control_conv2d_4 <= control_conv2d_4_11;
        end
        control_conv2d_4_11: begin
          if(cparam_conv2d_4_data_stationary == 0) begin
            control_conv2d_4 <= control_conv2d_4_12;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            control_conv2d_4 <= control_conv2d_4_24;
          end 
        end
        control_conv2d_4_12: begin
          control_conv2d_4 <= control_conv2d_4_13;
          if(conv2d_4_skip_read_act) begin
            control_conv2d_4 <= control_conv2d_4_23;
          end 
        end
        control_conv2d_4_13: begin
          control_conv2d_4 <= control_conv2d_4_14;
          if(conv2d_4_mux_dma_pad_mask_0 || !conv2d_4_mux_dma_flag_0) begin
            control_conv2d_4 <= control_conv2d_4_16;
          end 
        end
        control_conv2d_4_14: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_15;
          end 
        end
        control_conv2d_4_15: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_16;
          end 
        end
        control_conv2d_4_16: begin
          control_conv2d_4 <= control_conv2d_4_17;
          if(conv2d_4_mux_dma_pad_mask_1 || !conv2d_4_mux_dma_flag_1) begin
            control_conv2d_4 <= control_conv2d_4_19;
          end 
        end
        control_conv2d_4_17: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_18;
          end 
        end
        control_conv2d_4_18: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_19;
          end 
        end
        control_conv2d_4_19: begin
          control_conv2d_4 <= control_conv2d_4_20;
          if(conv2d_4_mux_dma_pad_mask_2 || !conv2d_4_mux_dma_flag_2) begin
            control_conv2d_4 <= control_conv2d_4_22;
          end 
        end
        control_conv2d_4_20: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_21;
          end 
        end
        control_conv2d_4_21: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_22;
          end 
        end
        control_conv2d_4_22: begin
          control_conv2d_4 <= control_conv2d_4_23;
        end
        control_conv2d_4_23: begin
          if(cparam_conv2d_4_data_stationary == 0) begin
            control_conv2d_4 <= control_conv2d_4_24;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            control_conv2d_4 <= control_conv2d_4_7;
          end 
        end
        control_conv2d_4_24: begin
          if(_maxi_write_idle) begin
            control_conv2d_4 <= control_conv2d_4_25;
          end 
        end
        control_conv2d_4_25: begin
          if(conv2d_4_comp_fsm == 0) begin
            control_conv2d_4 <= control_conv2d_4_26;
          end 
        end
        control_conv2d_4_26: begin
          control_conv2d_4 <= control_conv2d_4_27;
          if(conv2d_4_skip_write_out) begin
            control_conv2d_4 <= control_conv2d_4_32;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_prev_och_count < cparam_conv2d_4_max_och_count)) begin
            control_conv2d_4 <= control_conv2d_4_32;
          end 
        end
        control_conv2d_4_27: begin
          if(conv2d_4_sync_comp_count >= conv2d_4_sync_out_count + cparam_conv2d_4_inc_sync_out) begin
            control_conv2d_4 <= control_conv2d_4_28;
          end 
        end
        control_conv2d_4_28: begin
          if(!conv2d_4_dma_out_mask_0) begin
            control_conv2d_4 <= control_conv2d_4_29;
          end 
          if(conv2d_4_dma_out_mask_0) begin
            control_conv2d_4 <= control_conv2d_4_30;
          end 
        end
        control_conv2d_4_29: begin
          if(_maxi_write_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_30;
          end 
        end
        control_conv2d_4_30: begin
          control_conv2d_4 <= control_conv2d_4_31;
        end
        control_conv2d_4_31: begin
          conv2d_4_write_count <= conv2d_4_write_count + 1;
          if(conv2d_4_out_ram_select == 0) begin
            conv2d_4_out_laddr_offset <= conv2d_4_out_laddr_offset + conv2d_4_next_out_write_size;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !cparam_conv2d_4_keep_filter) begin
            conv2d_4_out_base_offset_col <= conv2d_4_out_base_offset_col + cparam_conv2d_4_out_col_step;
            conv2d_4_out_col_count <= conv2d_4_out_col_count + 1;
          end 
          conv2d_4_out_ram_select <= conv2d_4_out_ram_select + 1;
          if(conv2d_4_out_ram_select == 0) begin
            conv2d_4_out_ram_select <= 0;
          end 
          conv2d_4_sync_out_count <= conv2d_4_sync_out_count + cparam_conv2d_4_inc_sync_out;
          if((cparam_conv2d_4_data_stationary == 0) && !cparam_conv2d_4_keep_filter && (conv2d_4_write_count >= cparam_conv2d_4_out_num_col - 1) || (cparam_conv2d_4_data_stationary == 0) && cparam_conv2d_4_keep_filter || (cparam_conv2d_4_data_stationary == 1)) begin
            conv2d_4_sync_out_count <= conv2d_4_sync_out_count + (cparam_conv2d_4_inc_sync_out + cparam_conv2d_4_inc_sync_out_res);
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !cparam_conv2d_4_keep_filter) begin
            control_conv2d_4 <= control_conv2d_4_26;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !cparam_conv2d_4_keep_filter && (conv2d_4_write_count >= cparam_conv2d_4_out_num_col - 1) || (cparam_conv2d_4_data_stationary == 0) && cparam_conv2d_4_keep_filter || (cparam_conv2d_4_data_stationary == 1)) begin
            control_conv2d_4 <= control_conv2d_4_32;
          end 
        end
        control_conv2d_4_32: begin
          if(conv2d_4_update_filter) begin
            conv2d_4_filter_base_offset <= conv2d_4_filter_base_offset + cparam_conv2d_4_filter_base_step;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_filter_base_offset <= 0;
          end 
          if(conv2d_4_update_filter) begin
            conv2d_4_och_count <= conv2d_4_och_count + cparam_conv2d_4_och_count_step;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_och_count <= 0;
          end 
          if(conv2d_4_update_filter) begin
            conv2d_4_filter_page_comp_offset <= conv2d_4_filter_page_comp_offset + cparam_conv2d_4_filter_read_step;
            conv2d_4_filter_page_dma_offset <= conv2d_4_filter_page_dma_offset + cparam_conv2d_4_filter_read_step;
          end 
          if(conv2d_4_update_filter && (conv2d_4_filter_page_comp_offset + cparam_conv2d_4_filter_read_step + cparam_conv2d_4_filter_read_step > 512)) begin
            conv2d_4_filter_page_comp_offset <= 0;
            conv2d_4_filter_page_dma_offset <= 0;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_act_base_offset_row <= conv2d_4_act_base_offset_row + cparam_conv2d_4_act_row_step;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_act_base_offset_row <= 0;
            conv2d_4_act_base_offset_bat <= conv2d_4_act_base_offset_bat + cparam_conv2d_4_act_bat_step;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            conv2d_4_act_base_offset_bat <= 0;
          end 
          if(!conv2d_4_update_act) begin
            conv2d_4_dma_flag_0 <= 0;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_dma_flag_0 <= cparam_conv2d_4_dma_flag_conds_0;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_dma_flag_0 <= 1;
          end 
          if(!conv2d_4_update_act) begin
            conv2d_4_dma_flag_1 <= 0;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_dma_flag_1 <= cparam_conv2d_4_dma_flag_conds_1;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_dma_flag_1 <= 1;
          end 
          if(!conv2d_4_update_act) begin
            conv2d_4_dma_flag_2 <= 0;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_dma_flag_2 <= cparam_conv2d_4_dma_flag_conds_2;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_dma_flag_2 <= 1;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_row_count <= conv2d_4_row_count + cparam_conv2d_4_stride_row_par_row;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_row_count <= 0;
            conv2d_4_bat_count <= conv2d_4_bat_count + 1;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            conv2d_4_bat_count <= 0;
          end 
          if(conv2d_4_update_act && (cparam_conv2d_4_stride_row_par_row < 3)) begin
            conv2d_4_row_select <= conv2d_4_row_select + cparam_conv2d_4_stride_row_par_row;
            conv2d_4_prev_row_select <= conv2d_4_row_select;
          end 
          if(conv2d_4_update_act && (cparam_conv2d_4_stride_row_par_row < 3) && (conv2d_4_row_select + cparam_conv2d_4_stride_row_par_row >= 3)) begin
            conv2d_4_row_select <= conv2d_4_row_select - (3 - cparam_conv2d_4_stride_row_par_row);
            conv2d_4_prev_row_select <= conv2d_4_row_select;
          end 
          if(conv2d_4_update_act && !(cparam_conv2d_4_stride_row_par_row < 3)) begin
            conv2d_4_row_select <= 0;
            conv2d_4_prev_row_select <= 0;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_row_select <= 0;
            conv2d_4_prev_row_select <= 0;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_0) begin
            conv2d_4_act_page_comp_offset_0 <= conv2d_4_act_page_comp_offset_0 + cparam_conv2d_4_act_read_step;
            conv2d_4_act_page_dma_offset_0 <= conv2d_4_act_page_dma_offset_0 + cparam_conv2d_4_act_read_step;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_0 && (conv2d_4_act_page_comp_offset_0 + cparam_conv2d_4_act_read_step + cparam_conv2d_4_act_read_step > 1024)) begin
            conv2d_4_act_page_comp_offset_0 <= 0;
            conv2d_4_act_page_dma_offset_0 <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && cparam_conv2d_4_keep_input) begin
            conv2d_4_act_page_comp_offset_0 <= 0;
            conv2d_4_act_page_dma_offset_0 <= 0;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_1) begin
            conv2d_4_act_page_comp_offset_1 <= conv2d_4_act_page_comp_offset_1 + cparam_conv2d_4_act_read_step;
            conv2d_4_act_page_dma_offset_1 <= conv2d_4_act_page_dma_offset_1 + cparam_conv2d_4_act_read_step;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_1 && (conv2d_4_act_page_comp_offset_1 + cparam_conv2d_4_act_read_step + cparam_conv2d_4_act_read_step > 1024)) begin
            conv2d_4_act_page_comp_offset_1 <= 0;
            conv2d_4_act_page_dma_offset_1 <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && cparam_conv2d_4_keep_input) begin
            conv2d_4_act_page_comp_offset_1 <= 0;
            conv2d_4_act_page_dma_offset_1 <= 0;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_2) begin
            conv2d_4_act_page_comp_offset_2 <= conv2d_4_act_page_comp_offset_2 + cparam_conv2d_4_act_read_step;
            conv2d_4_act_page_dma_offset_2 <= conv2d_4_act_page_dma_offset_2 + cparam_conv2d_4_act_read_step;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_2 && (conv2d_4_act_page_comp_offset_2 + cparam_conv2d_4_act_read_step + cparam_conv2d_4_act_read_step > 1024)) begin
            conv2d_4_act_page_comp_offset_2 <= 0;
            conv2d_4_act_page_dma_offset_2 <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && cparam_conv2d_4_keep_input) begin
            conv2d_4_act_page_comp_offset_2 <= 0;
            conv2d_4_act_page_dma_offset_2 <= 0;
          end 
          conv2d_4_next_out_write_size <= (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)? cparam_conv2d_4_out_write_size_res : cparam_conv2d_4_out_write_size;
          if(!conv2d_4_skip_write_out) begin
            conv2d_4_write_count <= 0;
            conv2d_4_out_laddr_offset <= 0;
            conv2d_4_out_ram_select <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !conv2d_4_skip_write_out) begin
            conv2d_4_out_base_offset_col <= 0;
            conv2d_4_out_base_offset_row <= conv2d_4_out_base_offset_row + cparam_conv2d_4_out_row_step;
            conv2d_4_out_col_count <= 0;
            conv2d_4_out_row_count <= conv2d_4_out_row_count + 1;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !conv2d_4_skip_write_out && (conv2d_4_prev_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_out_base_offset_row <= 0;
            conv2d_4_out_base_offset_bat <= conv2d_4_out_base_offset_bat + cparam_conv2d_4_out_bat_step;
            conv2d_4_out_row_count <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !conv2d_4_skip_write_out && (conv2d_4_prev_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_prev_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            conv2d_4_out_base_offset_bat <= 0;
            conv2d_4_out_base_offset_och <= conv2d_4_out_base_offset_och + cparam_conv2d_4_out_och_step;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_prev_och_count >= cparam_conv2d_4_max_och_count) && !conv2d_4_skip_write_out) begin
            conv2d_4_out_base_offset_row <= conv2d_4_out_base_offset_row + cparam_conv2d_4_out_row_step;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !conv2d_4_out_page) begin
            conv2d_4_out_page_comp_offset <= 256;
            conv2d_4_out_page_dma_offset <= 0;
            conv2d_4_out_page <= 1;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && conv2d_4_out_page) begin
            conv2d_4_out_page_comp_offset <= 0;
            conv2d_4_out_page_dma_offset <= 256;
            conv2d_4_out_page <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count) && !conv2d_4_out_page) begin
            conv2d_4_out_page_comp_offset <= 256;
            conv2d_4_out_page_dma_offset <= 0;
            conv2d_4_out_page <= 1;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count) && conv2d_4_out_page) begin
            conv2d_4_out_page_comp_offset <= 0;
            conv2d_4_out_page_dma_offset <= 256;
            conv2d_4_out_page <= 0;
          end 
          conv2d_4_prev_row_count <= conv2d_4_row_count;
          conv2d_4_prev_bat_count <= conv2d_4_bat_count;
          conv2d_4_prev_och_count <= conv2d_4_och_count;
          if((conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_skip_read_filter <= 1;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && cparam_conv2d_4_keep_filter) begin
            conv2d_4_skip_read_filter <= 1;
          end 
          if((conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_skip_read_act <= 1;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && cparam_conv2d_4_keep_input) begin
            conv2d_4_skip_read_act <= 1;
          end 
          if((conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_skip_comp <= 1;
          end 
          if(conv2d_4_skip_write_out && (conv2d_4_prev_row_count == 0) && (conv2d_4_prev_bat_count == 0) && (conv2d_4_prev_och_count == 0)) begin
            conv2d_4_skip_write_out <= 0;
          end 
          if(cparam_conv2d_4_data_stationary == 0) begin
            control_conv2d_4 <= control_conv2d_4_12;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            control_conv2d_4 <= control_conv2d_4_7;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            control_conv2d_4 <= control_conv2d_4_7;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            control_conv2d_4 <= control_conv2d_4_12;
          end 
          if(!conv2d_4_skip_write_out && (conv2d_4_prev_och_count >= cparam_conv2d_4_max_och_count) && (conv2d_4_prev_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_prev_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            control_conv2d_4 <= control_conv2d_4_33;
          end 
        end
        control_conv2d_4_33: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_conv2d_4 <= control_conv2d_4_34;
          end 
        end
        control_conv2d_4_34: begin
          if(main_fsm == 14) begin
            _control_conv2d_4_called <= 0;
          end 
          if(main_fsm == 31) begin
            _control_conv2d_4_called <= 0;
          end 
          if(main_fsm == 48) begin
            _control_conv2d_4_called <= 0;
          end 
          if(main_fsm == 14) begin
            control_conv2d_4 <= control_conv2d_4_init;
          end 
          if(main_fsm == 31) begin
            control_conv2d_4 <= control_conv2d_4_init;
          end 
          if(main_fsm == 48) begin
            control_conv2d_4 <= control_conv2d_4_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_read_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_req_fsm <= _maxi_read_req_fsm_init;
      _maxi_read_cont <= 0;
    end else begin
      case(_maxi_read_req_fsm)
        _maxi_read_req_fsm_init: begin
          if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full) begin
            _maxi_read_req_fsm <= _maxi_read_req_fsm_1;
          end 
        end
        _maxi_read_req_fsm_1: begin
          if(maxi_arready || !maxi_arvalid) begin
            _maxi_read_cont <= 1;
          end 
          if((maxi_arready || !maxi_arvalid) && (_maxi_read_global_size == 0)) begin
            _maxi_read_cont <= 0;
          end 
          if(maxi_arready || !maxi_arvalid) begin
            _maxi_read_req_fsm <= _maxi_read_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_read_data_fsm_1 = 1;
  localparam _maxi_read_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
    end else begin
      case(_maxi_read_data_fsm)
        _maxi_read_data_fsm_init: begin
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 10)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 11)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 12)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 13)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 14)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 15)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
        end
        _maxi_read_data_fsm_1: begin
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
        end
        _maxi_read_data_fsm_2: begin
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_0_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_0 <= write_burst_packed_fsm_0_init;
      write_burst_packed_addr_79 <= 0;
      write_burst_packed_stride_80 <= 0;
      write_burst_packed_length_81 <= 0;
      write_burst_packed_done_82 <= 0;
    end else begin
      case(write_burst_packed_fsm_0)
        write_burst_packed_fsm_0_init: begin
          write_burst_packed_addr_79 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_80 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_81 <= _maxi_read_local_size_buf;
          write_burst_packed_done_82 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_0 <= write_burst_packed_fsm_0_1;
          end 
        end
        write_burst_packed_fsm_0_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_79 <= write_burst_packed_addr_79 + write_burst_packed_stride_80;
            write_burst_packed_length_81 <= write_burst_packed_length_81 - 1;
            write_burst_packed_done_82 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_81 <= 1)) begin
            write_burst_packed_done_82 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_82 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_81 <= 1)) begin
            write_burst_packed_fsm_0 <= write_burst_packed_fsm_0_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_0 <= write_burst_packed_fsm_0_init;
          end 
          if(0) begin
            write_burst_packed_fsm_0 <= write_burst_packed_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_1_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_init;
      write_burst_packed_addr_92 <= 0;
      write_burst_packed_stride_93 <= 0;
      write_burst_packed_length_94 <= 0;
      write_burst_packed_done_95 <= 0;
    end else begin
      case(write_burst_packed_fsm_1)
        write_burst_packed_fsm_1_init: begin
          write_burst_packed_addr_92 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_93 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_94 <= _maxi_read_local_size_buf;
          write_burst_packed_done_95 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 2) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_1;
          end 
        end
        write_burst_packed_fsm_1_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_92 <= write_burst_packed_addr_92 + write_burst_packed_stride_93;
            write_burst_packed_length_94 <= write_burst_packed_length_94 - 1;
            write_burst_packed_done_95 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_94 <= 1)) begin
            write_burst_packed_done_95 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_95 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_94 <= 1)) begin
            write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_init;
          end 
          if(0) begin
            write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_2_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_2 <= write_burst_packed_fsm_2_init;
      write_burst_packed_addr_110 <= 0;
      write_burst_packed_stride_111 <= 0;
      write_burst_packed_length_112 <= 0;
      write_burst_packed_done_113 <= 0;
    end else begin
      case(write_burst_packed_fsm_2)
        write_burst_packed_fsm_2_init: begin
          write_burst_packed_addr_110 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_111 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_112 <= _maxi_read_local_size_buf;
          write_burst_packed_done_113 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_2 <= write_burst_packed_fsm_2_1;
          end 
        end
        write_burst_packed_fsm_2_1: begin
          if(write_burst_block_ram_wvalid_108) begin
            write_burst_packed_addr_110 <= write_burst_packed_addr_110 + write_burst_packed_stride_111;
            write_burst_packed_length_112 <= write_burst_packed_length_112 - 1;
            write_burst_packed_done_113 <= 0;
          end 
          if(write_burst_block_ram_wvalid_108 && (write_burst_packed_length_112 <= 1)) begin
            write_burst_packed_done_113 <= 1;
          end 
          if(write_burst_block_ram_wvalid_108 && 0) begin
            write_burst_packed_done_113 <= 1;
          end 
          if(write_burst_block_ram_wvalid_108 && (write_burst_packed_length_112 <= 1)) begin
            write_burst_packed_fsm_2 <= write_burst_packed_fsm_2_init;
          end 
          if(write_burst_block_ram_wvalid_108 && 0) begin
            write_burst_packed_fsm_2 <= write_burst_packed_fsm_2_init;
          end 
          if(write_burst_block_ram_wquit_109) begin
            write_burst_packed_fsm_2 <= write_burst_packed_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_3_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_3 <= write_burst_packed_fsm_3_init;
      write_burst_packed_addr_120 <= 0;
      write_burst_packed_stride_121 <= 0;
      write_burst_packed_length_122 <= 0;
      write_burst_packed_done_123 <= 0;
    end else begin
      case(write_burst_packed_fsm_3)
        write_burst_packed_fsm_3_init: begin
          write_burst_packed_addr_120 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_121 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_122 <= _maxi_read_local_size_buf;
          write_burst_packed_done_123 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_3 <= write_burst_packed_fsm_3_1;
          end 
        end
        write_burst_packed_fsm_3_1: begin
          if(write_burst_block_ram_wvalid_118) begin
            write_burst_packed_addr_120 <= write_burst_packed_addr_120 + write_burst_packed_stride_121;
            write_burst_packed_length_122 <= write_burst_packed_length_122 - 1;
            write_burst_packed_done_123 <= 0;
          end 
          if(write_burst_block_ram_wvalid_118 && (write_burst_packed_length_122 <= 1)) begin
            write_burst_packed_done_123 <= 1;
          end 
          if(write_burst_block_ram_wvalid_118 && 0) begin
            write_burst_packed_done_123 <= 1;
          end 
          if(write_burst_block_ram_wvalid_118 && (write_burst_packed_length_122 <= 1)) begin
            write_burst_packed_fsm_3 <= write_burst_packed_fsm_3_init;
          end 
          if(write_burst_block_ram_wvalid_118 && 0) begin
            write_burst_packed_fsm_3 <= write_burst_packed_fsm_3_init;
          end 
          if(write_burst_block_ram_wquit_119) begin
            write_burst_packed_fsm_3 <= write_burst_packed_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_4_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_4 <= write_burst_packed_fsm_4_init;
      write_burst_packed_addr_130 <= 0;
      write_burst_packed_stride_131 <= 0;
      write_burst_packed_length_132 <= 0;
      write_burst_packed_done_133 <= 0;
    end else begin
      case(write_burst_packed_fsm_4)
        write_burst_packed_fsm_4_init: begin
          write_burst_packed_addr_130 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_131 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_132 <= _maxi_read_local_size_buf;
          write_burst_packed_done_133 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_4 <= write_burst_packed_fsm_4_1;
          end 
        end
        write_burst_packed_fsm_4_1: begin
          if(write_burst_block_ram_wvalid_128) begin
            write_burst_packed_addr_130 <= write_burst_packed_addr_130 + write_burst_packed_stride_131;
            write_burst_packed_length_132 <= write_burst_packed_length_132 - 1;
            write_burst_packed_done_133 <= 0;
          end 
          if(write_burst_block_ram_wvalid_128 && (write_burst_packed_length_132 <= 1)) begin
            write_burst_packed_done_133 <= 1;
          end 
          if(write_burst_block_ram_wvalid_128 && 0) begin
            write_burst_packed_done_133 <= 1;
          end 
          if(write_burst_block_ram_wvalid_128 && (write_burst_packed_length_132 <= 1)) begin
            write_burst_packed_fsm_4 <= write_burst_packed_fsm_4_init;
          end 
          if(write_burst_block_ram_wvalid_128 && 0) begin
            write_burst_packed_fsm_4 <= write_burst_packed_fsm_4_init;
          end 
          if(write_burst_block_ram_wquit_129) begin
            write_burst_packed_fsm_4 <= write_burst_packed_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_5_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_init;
      write_burst_packed_addr_140 <= 0;
      write_burst_packed_stride_141 <= 0;
      write_burst_packed_length_142 <= 0;
      write_burst_packed_done_143 <= 0;
    end else begin
      case(write_burst_packed_fsm_5)
        write_burst_packed_fsm_5_init: begin
          write_burst_packed_addr_140 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_141 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_142 <= _maxi_read_local_size_buf;
          write_burst_packed_done_143 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_1;
          end 
        end
        write_burst_packed_fsm_5_1: begin
          if(write_burst_block_ram_wvalid_138) begin
            write_burst_packed_addr_140 <= write_burst_packed_addr_140 + write_burst_packed_stride_141;
            write_burst_packed_length_142 <= write_burst_packed_length_142 - 1;
            write_burst_packed_done_143 <= 0;
          end 
          if(write_burst_block_ram_wvalid_138 && (write_burst_packed_length_142 <= 1)) begin
            write_burst_packed_done_143 <= 1;
          end 
          if(write_burst_block_ram_wvalid_138 && 0) begin
            write_burst_packed_done_143 <= 1;
          end 
          if(write_burst_block_ram_wvalid_138 && (write_burst_packed_length_142 <= 1)) begin
            write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_init;
          end 
          if(write_burst_block_ram_wvalid_138 && 0) begin
            write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_init;
          end 
          if(write_burst_block_ram_wquit_139) begin
            write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_6_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_6 <= write_burst_packed_fsm_6_init;
      write_burst_packed_addr_150 <= 0;
      write_burst_packed_stride_151 <= 0;
      write_burst_packed_length_152 <= 0;
      write_burst_packed_done_153 <= 0;
    end else begin
      case(write_burst_packed_fsm_6)
        write_burst_packed_fsm_6_init: begin
          write_burst_packed_addr_150 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_151 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_152 <= _maxi_read_local_size_buf;
          write_burst_packed_done_153 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_6 <= write_burst_packed_fsm_6_1;
          end 
        end
        write_burst_packed_fsm_6_1: begin
          if(write_burst_block_ram_wvalid_148) begin
            write_burst_packed_addr_150 <= write_burst_packed_addr_150 + write_burst_packed_stride_151;
            write_burst_packed_length_152 <= write_burst_packed_length_152 - 1;
            write_burst_packed_done_153 <= 0;
          end 
          if(write_burst_block_ram_wvalid_148 && (write_burst_packed_length_152 <= 1)) begin
            write_burst_packed_done_153 <= 1;
          end 
          if(write_burst_block_ram_wvalid_148 && 0) begin
            write_burst_packed_done_153 <= 1;
          end 
          if(write_burst_block_ram_wvalid_148 && (write_burst_packed_length_152 <= 1)) begin
            write_burst_packed_fsm_6 <= write_burst_packed_fsm_6_init;
          end 
          if(write_burst_block_ram_wvalid_148 && 0) begin
            write_burst_packed_fsm_6 <= write_burst_packed_fsm_6_init;
          end 
          if(write_burst_block_ram_wquit_149) begin
            write_burst_packed_fsm_6 <= write_burst_packed_fsm_6_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_7_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_7 <= write_burst_packed_fsm_7_init;
      write_burst_packed_addr_160 <= 0;
      write_burst_packed_stride_161 <= 0;
      write_burst_packed_length_162 <= 0;
      write_burst_packed_done_163 <= 0;
    end else begin
      case(write_burst_packed_fsm_7)
        write_burst_packed_fsm_7_init: begin
          write_burst_packed_addr_160 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_161 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_162 <= _maxi_read_local_size_buf;
          write_burst_packed_done_163 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_7 <= write_burst_packed_fsm_7_1;
          end 
        end
        write_burst_packed_fsm_7_1: begin
          if(write_burst_block_ram_wvalid_158) begin
            write_burst_packed_addr_160 <= write_burst_packed_addr_160 + write_burst_packed_stride_161;
            write_burst_packed_length_162 <= write_burst_packed_length_162 - 1;
            write_burst_packed_done_163 <= 0;
          end 
          if(write_burst_block_ram_wvalid_158 && (write_burst_packed_length_162 <= 1)) begin
            write_burst_packed_done_163 <= 1;
          end 
          if(write_burst_block_ram_wvalid_158 && 0) begin
            write_burst_packed_done_163 <= 1;
          end 
          if(write_burst_block_ram_wvalid_158 && (write_burst_packed_length_162 <= 1)) begin
            write_burst_packed_fsm_7 <= write_burst_packed_fsm_7_init;
          end 
          if(write_burst_block_ram_wvalid_158 && 0) begin
            write_burst_packed_fsm_7 <= write_burst_packed_fsm_7_init;
          end 
          if(write_burst_block_ram_wquit_159) begin
            write_burst_packed_fsm_7 <= write_burst_packed_fsm_7_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_8_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_8 <= write_burst_packed_fsm_8_init;
      write_burst_packed_addr_170 <= 0;
      write_burst_packed_stride_171 <= 0;
      write_burst_packed_length_172 <= 0;
      write_burst_packed_done_173 <= 0;
    end else begin
      case(write_burst_packed_fsm_8)
        write_burst_packed_fsm_8_init: begin
          write_burst_packed_addr_170 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_171 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_172 <= _maxi_read_local_size_buf;
          write_burst_packed_done_173 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_8 <= write_burst_packed_fsm_8_1;
          end 
        end
        write_burst_packed_fsm_8_1: begin
          if(write_burst_block_ram_wvalid_168) begin
            write_burst_packed_addr_170 <= write_burst_packed_addr_170 + write_burst_packed_stride_171;
            write_burst_packed_length_172 <= write_burst_packed_length_172 - 1;
            write_burst_packed_done_173 <= 0;
          end 
          if(write_burst_block_ram_wvalid_168 && (write_burst_packed_length_172 <= 1)) begin
            write_burst_packed_done_173 <= 1;
          end 
          if(write_burst_block_ram_wvalid_168 && 0) begin
            write_burst_packed_done_173 <= 1;
          end 
          if(write_burst_block_ram_wvalid_168 && (write_burst_packed_length_172 <= 1)) begin
            write_burst_packed_fsm_8 <= write_burst_packed_fsm_8_init;
          end 
          if(write_burst_block_ram_wvalid_168 && 0) begin
            write_burst_packed_fsm_8 <= write_burst_packed_fsm_8_init;
          end 
          if(write_burst_block_ram_wquit_169) begin
            write_burst_packed_fsm_8 <= write_burst_packed_fsm_8_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_9_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_9 <= write_burst_packed_fsm_9_init;
      write_burst_packed_addr_180 <= 0;
      write_burst_packed_stride_181 <= 0;
      write_burst_packed_length_182 <= 0;
      write_burst_packed_done_183 <= 0;
    end else begin
      case(write_burst_packed_fsm_9)
        write_burst_packed_fsm_9_init: begin
          write_burst_packed_addr_180 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_181 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_182 <= _maxi_read_local_size_buf;
          write_burst_packed_done_183 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_9 <= write_burst_packed_fsm_9_1;
          end 
        end
        write_burst_packed_fsm_9_1: begin
          if(write_burst_block_ram_wvalid_178) begin
            write_burst_packed_addr_180 <= write_burst_packed_addr_180 + write_burst_packed_stride_181;
            write_burst_packed_length_182 <= write_burst_packed_length_182 - 1;
            write_burst_packed_done_183 <= 0;
          end 
          if(write_burst_block_ram_wvalid_178 && (write_burst_packed_length_182 <= 1)) begin
            write_burst_packed_done_183 <= 1;
          end 
          if(write_burst_block_ram_wvalid_178 && 0) begin
            write_burst_packed_done_183 <= 1;
          end 
          if(write_burst_block_ram_wvalid_178 && (write_burst_packed_length_182 <= 1)) begin
            write_burst_packed_fsm_9 <= write_burst_packed_fsm_9_init;
          end 
          if(write_burst_block_ram_wvalid_178 && 0) begin
            write_burst_packed_fsm_9 <= write_burst_packed_fsm_9_init;
          end 
          if(write_burst_block_ram_wquit_179) begin
            write_burst_packed_fsm_9 <= write_burst_packed_fsm_9_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_10_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_10 <= write_burst_packed_fsm_10_init;
      write_burst_packed_addr_190 <= 0;
      write_burst_packed_stride_191 <= 0;
      write_burst_packed_length_192 <= 0;
      write_burst_packed_done_193 <= 0;
    end else begin
      case(write_burst_packed_fsm_10)
        write_burst_packed_fsm_10_init: begin
          write_burst_packed_addr_190 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_191 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_192 <= _maxi_read_local_size_buf;
          write_burst_packed_done_193 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_10 <= write_burst_packed_fsm_10_1;
          end 
        end
        write_burst_packed_fsm_10_1: begin
          if(write_burst_block_ram_wvalid_188) begin
            write_burst_packed_addr_190 <= write_burst_packed_addr_190 + write_burst_packed_stride_191;
            write_burst_packed_length_192 <= write_burst_packed_length_192 - 1;
            write_burst_packed_done_193 <= 0;
          end 
          if(write_burst_block_ram_wvalid_188 && (write_burst_packed_length_192 <= 1)) begin
            write_burst_packed_done_193 <= 1;
          end 
          if(write_burst_block_ram_wvalid_188 && 0) begin
            write_burst_packed_done_193 <= 1;
          end 
          if(write_burst_block_ram_wvalid_188 && (write_burst_packed_length_192 <= 1)) begin
            write_burst_packed_fsm_10 <= write_burst_packed_fsm_10_init;
          end 
          if(write_burst_block_ram_wvalid_188 && 0) begin
            write_burst_packed_fsm_10 <= write_burst_packed_fsm_10_init;
          end 
          if(write_burst_block_ram_wquit_189) begin
            write_burst_packed_fsm_10 <= write_burst_packed_fsm_10_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_11_1 = 1;
  localparam write_burst_block_fsm_11_2 = 2;
  localparam write_burst_block_fsm_11_3 = 3;
  localparam write_burst_block_fsm_11_4 = 4;
  localparam write_burst_block_fsm_11_5 = 5;
  localparam write_burst_block_fsm_11_6 = 6;
  localparam write_burst_block_fsm_11_7 = 7;
  localparam write_burst_block_fsm_11_8 = 8;
  localparam write_burst_block_fsm_11_9 = 9;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
      write_burst_block_length_198 <= 0;
      write_burst_block_blocksize_199 <= 0;
      write_burst_block_done_200 <= 0;
      write_burst_block_count_201 <= 0;
    end else begin
      case(write_burst_block_fsm_11)
        write_burst_block_fsm_11_init: begin
          write_burst_block_length_198 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_199 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_200 <= 0;
          write_burst_block_count_201 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_1;
          end 
        end
        write_burst_block_fsm_11_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_4;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_4: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_5;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_5: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_6;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_6: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_7;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_7: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_8;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_8: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_9;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_9: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_12_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_12 <= write_burst_packed_fsm_12_init;
      write_burst_packed_addr_212 <= 0;
      write_burst_packed_stride_213 <= 0;
      write_burst_packed_length_214 <= 0;
      write_burst_packed_done_215 <= 0;
    end else begin
      case(write_burst_packed_fsm_12)
        write_burst_packed_fsm_12_init: begin
          write_burst_packed_addr_212 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_213 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_214 <= _maxi_read_local_size_buf;
          write_burst_packed_done_215 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_12 <= write_burst_packed_fsm_12_1;
          end 
        end
        write_burst_packed_fsm_12_1: begin
          if(write_burst_block_ram_wvalid_210) begin
            write_burst_packed_addr_212 <= write_burst_packed_addr_212 + write_burst_packed_stride_213;
            write_burst_packed_length_214 <= write_burst_packed_length_214 - 1;
            write_burst_packed_done_215 <= 0;
          end 
          if(write_burst_block_ram_wvalid_210 && (write_burst_packed_length_214 <= 1)) begin
            write_burst_packed_done_215 <= 1;
          end 
          if(write_burst_block_ram_wvalid_210 && 0) begin
            write_burst_packed_done_215 <= 1;
          end 
          if(write_burst_block_ram_wvalid_210 && (write_burst_packed_length_214 <= 1)) begin
            write_burst_packed_fsm_12 <= write_burst_packed_fsm_12_init;
          end 
          if(write_burst_block_ram_wvalid_210 && 0) begin
            write_burst_packed_fsm_12 <= write_burst_packed_fsm_12_init;
          end 
          if(write_burst_block_ram_wquit_211) begin
            write_burst_packed_fsm_12 <= write_burst_packed_fsm_12_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_13_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_13 <= write_burst_packed_fsm_13_init;
      write_burst_packed_addr_222 <= 0;
      write_burst_packed_stride_223 <= 0;
      write_burst_packed_length_224 <= 0;
      write_burst_packed_done_225 <= 0;
    end else begin
      case(write_burst_packed_fsm_13)
        write_burst_packed_fsm_13_init: begin
          write_burst_packed_addr_222 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_223 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_224 <= _maxi_read_local_size_buf;
          write_burst_packed_done_225 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_13 <= write_burst_packed_fsm_13_1;
          end 
        end
        write_burst_packed_fsm_13_1: begin
          if(write_burst_block_ram_wvalid_220) begin
            write_burst_packed_addr_222 <= write_burst_packed_addr_222 + write_burst_packed_stride_223;
            write_burst_packed_length_224 <= write_burst_packed_length_224 - 1;
            write_burst_packed_done_225 <= 0;
          end 
          if(write_burst_block_ram_wvalid_220 && (write_burst_packed_length_224 <= 1)) begin
            write_burst_packed_done_225 <= 1;
          end 
          if(write_burst_block_ram_wvalid_220 && 0) begin
            write_burst_packed_done_225 <= 1;
          end 
          if(write_burst_block_ram_wvalid_220 && (write_burst_packed_length_224 <= 1)) begin
            write_burst_packed_fsm_13 <= write_burst_packed_fsm_13_init;
          end 
          if(write_burst_block_ram_wvalid_220 && 0) begin
            write_burst_packed_fsm_13 <= write_burst_packed_fsm_13_init;
          end 
          if(write_burst_block_ram_wquit_221) begin
            write_burst_packed_fsm_13 <= write_burst_packed_fsm_13_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_14_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_14 <= write_burst_packed_fsm_14_init;
      write_burst_packed_addr_232 <= 0;
      write_burst_packed_stride_233 <= 0;
      write_burst_packed_length_234 <= 0;
      write_burst_packed_done_235 <= 0;
    end else begin
      case(write_burst_packed_fsm_14)
        write_burst_packed_fsm_14_init: begin
          write_burst_packed_addr_232 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_233 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_234 <= _maxi_read_local_size_buf;
          write_burst_packed_done_235 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_14 <= write_burst_packed_fsm_14_1;
          end 
        end
        write_burst_packed_fsm_14_1: begin
          if(write_burst_block_ram_wvalid_230) begin
            write_burst_packed_addr_232 <= write_burst_packed_addr_232 + write_burst_packed_stride_233;
            write_burst_packed_length_234 <= write_burst_packed_length_234 - 1;
            write_burst_packed_done_235 <= 0;
          end 
          if(write_burst_block_ram_wvalid_230 && (write_burst_packed_length_234 <= 1)) begin
            write_burst_packed_done_235 <= 1;
          end 
          if(write_burst_block_ram_wvalid_230 && 0) begin
            write_burst_packed_done_235 <= 1;
          end 
          if(write_burst_block_ram_wvalid_230 && (write_burst_packed_length_234 <= 1)) begin
            write_burst_packed_fsm_14 <= write_burst_packed_fsm_14_init;
          end 
          if(write_burst_block_ram_wvalid_230 && 0) begin
            write_burst_packed_fsm_14 <= write_burst_packed_fsm_14_init;
          end 
          if(write_burst_block_ram_wquit_231) begin
            write_burst_packed_fsm_14 <= write_burst_packed_fsm_14_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_15_1 = 1;
  localparam write_burst_block_fsm_15_2 = 2;
  localparam write_burst_block_fsm_15_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
      write_burst_block_length_240 <= 0;
      write_burst_block_blocksize_241 <= 0;
      write_burst_block_done_242 <= 0;
      write_burst_block_count_243 <= 0;
    end else begin
      case(write_burst_block_fsm_15)
        write_burst_block_fsm_15_init: begin
          write_burst_block_length_240 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_241 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_242 <= 0;
          write_burst_block_count_243 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_1;
          end 
        end
        write_burst_block_fsm_15_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_240 <= write_burst_block_length_240 - 1;
            write_burst_block_done_242 <= 0;
            write_burst_block_count_243 <= write_burst_block_count_243 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1)) begin
            write_burst_block_done_242 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_242 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_243 == write_burst_block_blocksize_241 - 1)) begin
            write_burst_block_count_243 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_243 == write_burst_block_blocksize_241 - 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
        end
        write_burst_block_fsm_15_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_240 <= write_burst_block_length_240 - 1;
            write_burst_block_done_242 <= 0;
            write_burst_block_count_243 <= write_burst_block_count_243 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1)) begin
            write_burst_block_done_242 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_242 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_243 == write_burst_block_blocksize_241 - 1)) begin
            write_burst_block_count_243 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_243 == write_burst_block_blocksize_241 - 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
        end
        write_burst_block_fsm_15_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_240 <= write_burst_block_length_240 - 1;
            write_burst_block_done_242 <= 0;
            write_burst_block_count_243 <= write_burst_block_count_243 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1)) begin
            write_burst_block_done_242 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_242 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_243 == write_burst_block_blocksize_241 - 1)) begin
            write_burst_block_count_243 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_243 == write_burst_block_blocksize_241 - 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_16_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_16 <= write_burst_packed_fsm_16_init;
      write_burst_packed_addr_254 <= 0;
      write_burst_packed_stride_255 <= 0;
      write_burst_packed_length_256 <= 0;
      write_burst_packed_done_257 <= 0;
    end else begin
      case(write_burst_packed_fsm_16)
        write_burst_packed_fsm_16_init: begin
          write_burst_packed_addr_254 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_255 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_256 <= _maxi_read_local_size_buf;
          write_burst_packed_done_257 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_16 <= write_burst_packed_fsm_16_1;
          end 
        end
        write_burst_packed_fsm_16_1: begin
          if(write_burst_block_ram_wvalid_252) begin
            write_burst_packed_addr_254 <= write_burst_packed_addr_254 + write_burst_packed_stride_255;
            write_burst_packed_length_256 <= write_burst_packed_length_256 - 1;
            write_burst_packed_done_257 <= 0;
          end 
          if(write_burst_block_ram_wvalid_252 && (write_burst_packed_length_256 <= 1)) begin
            write_burst_packed_done_257 <= 1;
          end 
          if(write_burst_block_ram_wvalid_252 && 0) begin
            write_burst_packed_done_257 <= 1;
          end 
          if(write_burst_block_ram_wvalid_252 && (write_burst_packed_length_256 <= 1)) begin
            write_burst_packed_fsm_16 <= write_burst_packed_fsm_16_init;
          end 
          if(write_burst_block_ram_wvalid_252 && 0) begin
            write_burst_packed_fsm_16 <= write_burst_packed_fsm_16_init;
          end 
          if(write_burst_block_ram_wquit_253) begin
            write_burst_packed_fsm_16 <= write_burst_packed_fsm_16_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_17_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_17 <= write_burst_packed_fsm_17_init;
      write_burst_packed_addr_264 <= 0;
      write_burst_packed_stride_265 <= 0;
      write_burst_packed_length_266 <= 0;
      write_burst_packed_done_267 <= 0;
    end else begin
      case(write_burst_packed_fsm_17)
        write_burst_packed_fsm_17_init: begin
          write_burst_packed_addr_264 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_265 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_266 <= _maxi_read_local_size_buf;
          write_burst_packed_done_267 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_17 <= write_burst_packed_fsm_17_1;
          end 
        end
        write_burst_packed_fsm_17_1: begin
          if(write_burst_block_ram_wvalid_262) begin
            write_burst_packed_addr_264 <= write_burst_packed_addr_264 + write_burst_packed_stride_265;
            write_burst_packed_length_266 <= write_burst_packed_length_266 - 1;
            write_burst_packed_done_267 <= 0;
          end 
          if(write_burst_block_ram_wvalid_262 && (write_burst_packed_length_266 <= 1)) begin
            write_burst_packed_done_267 <= 1;
          end 
          if(write_burst_block_ram_wvalid_262 && 0) begin
            write_burst_packed_done_267 <= 1;
          end 
          if(write_burst_block_ram_wvalid_262 && (write_burst_packed_length_266 <= 1)) begin
            write_burst_packed_fsm_17 <= write_burst_packed_fsm_17_init;
          end 
          if(write_burst_block_ram_wvalid_262 && 0) begin
            write_burst_packed_fsm_17 <= write_burst_packed_fsm_17_init;
          end 
          if(write_burst_block_ram_wquit_263) begin
            write_burst_packed_fsm_17 <= write_burst_packed_fsm_17_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_18_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_18 <= write_burst_packed_fsm_18_init;
      write_burst_packed_addr_274 <= 0;
      write_burst_packed_stride_275 <= 0;
      write_burst_packed_length_276 <= 0;
      write_burst_packed_done_277 <= 0;
    end else begin
      case(write_burst_packed_fsm_18)
        write_burst_packed_fsm_18_init: begin
          write_burst_packed_addr_274 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_275 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_276 <= _maxi_read_local_size_buf;
          write_burst_packed_done_277 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_18 <= write_burst_packed_fsm_18_1;
          end 
        end
        write_burst_packed_fsm_18_1: begin
          if(write_burst_block_ram_wvalid_272) begin
            write_burst_packed_addr_274 <= write_burst_packed_addr_274 + write_burst_packed_stride_275;
            write_burst_packed_length_276 <= write_burst_packed_length_276 - 1;
            write_burst_packed_done_277 <= 0;
          end 
          if(write_burst_block_ram_wvalid_272 && (write_burst_packed_length_276 <= 1)) begin
            write_burst_packed_done_277 <= 1;
          end 
          if(write_burst_block_ram_wvalid_272 && 0) begin
            write_burst_packed_done_277 <= 1;
          end 
          if(write_burst_block_ram_wvalid_272 && (write_burst_packed_length_276 <= 1)) begin
            write_burst_packed_fsm_18 <= write_burst_packed_fsm_18_init;
          end 
          if(write_burst_block_ram_wvalid_272 && 0) begin
            write_burst_packed_fsm_18 <= write_burst_packed_fsm_18_init;
          end 
          if(write_burst_block_ram_wquit_273) begin
            write_burst_packed_fsm_18 <= write_burst_packed_fsm_18_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_19_1 = 1;
  localparam write_burst_block_fsm_19_2 = 2;
  localparam write_burst_block_fsm_19_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
      write_burst_block_length_282 <= 0;
      write_burst_block_blocksize_283 <= 0;
      write_burst_block_done_284 <= 0;
      write_burst_block_count_285 <= 0;
    end else begin
      case(write_burst_block_fsm_19)
        write_burst_block_fsm_19_init: begin
          write_burst_block_length_282 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_283 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_284 <= 0;
          write_burst_block_count_285 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_1;
          end 
        end
        write_burst_block_fsm_19_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_282 <= write_burst_block_length_282 - 1;
            write_burst_block_done_284 <= 0;
            write_burst_block_count_285 <= write_burst_block_count_285 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1)) begin
            write_burst_block_done_284 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_284 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_285 == write_burst_block_blocksize_283 - 1)) begin
            write_burst_block_count_285 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_285 == write_burst_block_blocksize_283 - 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
        end
        write_burst_block_fsm_19_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_282 <= write_burst_block_length_282 - 1;
            write_burst_block_done_284 <= 0;
            write_burst_block_count_285 <= write_burst_block_count_285 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1)) begin
            write_burst_block_done_284 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_284 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_285 == write_burst_block_blocksize_283 - 1)) begin
            write_burst_block_count_285 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_285 == write_burst_block_blocksize_283 - 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
        end
        write_burst_block_fsm_19_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_282 <= write_burst_block_length_282 - 1;
            write_burst_block_done_284 <= 0;
            write_burst_block_count_285 <= write_burst_block_count_285 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1)) begin
            write_burst_block_done_284 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_284 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_285 == write_burst_block_blocksize_283 - 1)) begin
            write_burst_block_count_285 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_285 == write_burst_block_blocksize_283 - 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_20_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_20 <= write_burst_packed_fsm_20_init;
      write_burst_packed_addr_296 <= 0;
      write_burst_packed_stride_297 <= 0;
      write_burst_packed_length_298 <= 0;
      write_burst_packed_done_299 <= 0;
    end else begin
      case(write_burst_packed_fsm_20)
        write_burst_packed_fsm_20_init: begin
          write_burst_packed_addr_296 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_297 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_298 <= _maxi_read_local_size_buf;
          write_burst_packed_done_299 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_20 <= write_burst_packed_fsm_20_1;
          end 
        end
        write_burst_packed_fsm_20_1: begin
          if(write_burst_block_ram_wvalid_294) begin
            write_burst_packed_addr_296 <= write_burst_packed_addr_296 + write_burst_packed_stride_297;
            write_burst_packed_length_298 <= write_burst_packed_length_298 - 1;
            write_burst_packed_done_299 <= 0;
          end 
          if(write_burst_block_ram_wvalid_294 && (write_burst_packed_length_298 <= 1)) begin
            write_burst_packed_done_299 <= 1;
          end 
          if(write_burst_block_ram_wvalid_294 && 0) begin
            write_burst_packed_done_299 <= 1;
          end 
          if(write_burst_block_ram_wvalid_294 && (write_burst_packed_length_298 <= 1)) begin
            write_burst_packed_fsm_20 <= write_burst_packed_fsm_20_init;
          end 
          if(write_burst_block_ram_wvalid_294 && 0) begin
            write_burst_packed_fsm_20 <= write_burst_packed_fsm_20_init;
          end 
          if(write_burst_block_ram_wquit_295) begin
            write_burst_packed_fsm_20 <= write_burst_packed_fsm_20_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_21_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_21 <= write_burst_packed_fsm_21_init;
      write_burst_packed_addr_306 <= 0;
      write_burst_packed_stride_307 <= 0;
      write_burst_packed_length_308 <= 0;
      write_burst_packed_done_309 <= 0;
    end else begin
      case(write_burst_packed_fsm_21)
        write_burst_packed_fsm_21_init: begin
          write_burst_packed_addr_306 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_307 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_308 <= _maxi_read_local_size_buf;
          write_burst_packed_done_309 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_21 <= write_burst_packed_fsm_21_1;
          end 
        end
        write_burst_packed_fsm_21_1: begin
          if(write_burst_block_ram_wvalid_304) begin
            write_burst_packed_addr_306 <= write_burst_packed_addr_306 + write_burst_packed_stride_307;
            write_burst_packed_length_308 <= write_burst_packed_length_308 - 1;
            write_burst_packed_done_309 <= 0;
          end 
          if(write_burst_block_ram_wvalid_304 && (write_burst_packed_length_308 <= 1)) begin
            write_burst_packed_done_309 <= 1;
          end 
          if(write_burst_block_ram_wvalid_304 && 0) begin
            write_burst_packed_done_309 <= 1;
          end 
          if(write_burst_block_ram_wvalid_304 && (write_burst_packed_length_308 <= 1)) begin
            write_burst_packed_fsm_21 <= write_burst_packed_fsm_21_init;
          end 
          if(write_burst_block_ram_wvalid_304 && 0) begin
            write_burst_packed_fsm_21 <= write_burst_packed_fsm_21_init;
          end 
          if(write_burst_block_ram_wquit_305) begin
            write_burst_packed_fsm_21 <= write_burst_packed_fsm_21_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_22_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_22 <= write_burst_packed_fsm_22_init;
      write_burst_packed_addr_316 <= 0;
      write_burst_packed_stride_317 <= 0;
      write_burst_packed_length_318 <= 0;
      write_burst_packed_done_319 <= 0;
    end else begin
      case(write_burst_packed_fsm_22)
        write_burst_packed_fsm_22_init: begin
          write_burst_packed_addr_316 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_317 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_318 <= _maxi_read_local_size_buf;
          write_burst_packed_done_319 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_22 <= write_burst_packed_fsm_22_1;
          end 
        end
        write_burst_packed_fsm_22_1: begin
          if(write_burst_block_ram_wvalid_314) begin
            write_burst_packed_addr_316 <= write_burst_packed_addr_316 + write_burst_packed_stride_317;
            write_burst_packed_length_318 <= write_burst_packed_length_318 - 1;
            write_burst_packed_done_319 <= 0;
          end 
          if(write_burst_block_ram_wvalid_314 && (write_burst_packed_length_318 <= 1)) begin
            write_burst_packed_done_319 <= 1;
          end 
          if(write_burst_block_ram_wvalid_314 && 0) begin
            write_burst_packed_done_319 <= 1;
          end 
          if(write_burst_block_ram_wvalid_314 && (write_burst_packed_length_318 <= 1)) begin
            write_burst_packed_fsm_22 <= write_burst_packed_fsm_22_init;
          end 
          if(write_burst_block_ram_wvalid_314 && 0) begin
            write_burst_packed_fsm_22 <= write_burst_packed_fsm_22_init;
          end 
          if(write_burst_block_ram_wquit_315) begin
            write_burst_packed_fsm_22 <= write_burst_packed_fsm_22_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_23_1 = 1;
  localparam write_burst_block_fsm_23_2 = 2;
  localparam write_burst_block_fsm_23_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
      write_burst_block_length_324 <= 0;
      write_burst_block_blocksize_325 <= 0;
      write_burst_block_done_326 <= 0;
      write_burst_block_count_327 <= 0;
    end else begin
      case(write_burst_block_fsm_23)
        write_burst_block_fsm_23_init: begin
          write_burst_block_length_324 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_325 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_326 <= 0;
          write_burst_block_count_327 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_1;
          end 
        end
        write_burst_block_fsm_23_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_324 <= write_burst_block_length_324 - 1;
            write_burst_block_done_326 <= 0;
            write_burst_block_count_327 <= write_burst_block_count_327 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1)) begin
            write_burst_block_done_326 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_326 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_327 == write_burst_block_blocksize_325 - 1)) begin
            write_burst_block_count_327 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_327 == write_burst_block_blocksize_325 - 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
        end
        write_burst_block_fsm_23_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_324 <= write_burst_block_length_324 - 1;
            write_burst_block_done_326 <= 0;
            write_burst_block_count_327 <= write_burst_block_count_327 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1)) begin
            write_burst_block_done_326 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_326 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_327 == write_burst_block_blocksize_325 - 1)) begin
            write_burst_block_count_327 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_327 == write_burst_block_blocksize_325 - 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
        end
        write_burst_block_fsm_23_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_324 <= write_burst_block_length_324 - 1;
            write_burst_block_done_326 <= 0;
            write_burst_block_count_327 <= write_burst_block_count_327 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1)) begin
            write_burst_block_done_326 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_326 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_327 == write_burst_block_blocksize_325 - 1)) begin
            write_burst_block_count_327 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_327 == write_burst_block_blocksize_325 - 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
        end
      endcase
    end
  end

  localparam conv2d_4_comp_fsm_1 = 1;
  localparam conv2d_4_comp_fsm_2 = 2;
  localparam conv2d_4_comp_fsm_3 = 3;
  localparam conv2d_4_comp_fsm_4 = 4;
  localparam conv2d_4_comp_fsm_5 = 5;
  localparam conv2d_4_comp_fsm_6 = 6;

  always @(posedge CLK) begin
    if(RST) begin
      conv2d_4_comp_fsm <= conv2d_4_comp_fsm_init;
      conv2d_4_stream_act_local_0 <= 0;
      conv2d_4_stream_act_local_1 <= 0;
      conv2d_4_stream_act_local_2 <= 0;
      conv2d_4_stream_act_local_3 <= 0;
      conv2d_4_stream_act_local_4 <= 0;
      conv2d_4_stream_act_local_5 <= 0;
      conv2d_4_stream_act_local_6 <= 0;
      conv2d_4_stream_act_local_7 <= 0;
      conv2d_4_stream_act_local_8 <= 0;
      conv2d_4_stream_out_local_col <= 0;
      conv2d_4_stream_out_local_val <= 0;
      conv2d_4_col_count <= 0;
      conv2d_4_col_select <= 0;
      conv2d_4_filter_page_comp_offset_buf <= 0;
      conv2d_4_act_page_comp_offset_buf_0 <= 0;
      conv2d_4_act_page_comp_offset_buf_1 <= 0;
      conv2d_4_act_page_comp_offset_buf_2 <= 0;
      conv2d_4_out_page_comp_offset_buf <= 0;
      conv2d_4_row_count_buf <= 0;
      conv2d_4_row_select_buf <= 0;
      conv2d_4_och_count_buf <= 0;
      conv2d_4_next_stream_num_ops <= 0;
      conv2d_4_stream_pad_masks <= 0;
      conv2d_4_sync_comp_count <= 0;
    end else begin
      if(_stream_conv2d_4_sink_stop) begin
        conv2d_4_sync_comp_count <= conv2d_4_sync_comp_count + 1;
      end 
      if(control_conv2d_4 == 6) begin
        conv2d_4_sync_comp_count <= 0;
      end 
      case(conv2d_4_comp_fsm)
        conv2d_4_comp_fsm_init: begin
          if((control_conv2d_4 == 25) && !conv2d_4_skip_comp) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_1;
          end 
        end
        conv2d_4_comp_fsm_1: begin
          conv2d_4_stream_act_local_0 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_0 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_0 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_1 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_1 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_1 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_2 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_2 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_2 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_3 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_3 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_3 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_4 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_4 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_4 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_5 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_5 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_5 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_6 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_6 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_6 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_7 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_7 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_7 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_8 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_8 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_8 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_out_local_col <= 0;
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count == 0)) begin
            conv2d_4_stream_out_local_val <= 0;
          end 
          conv2d_4_col_count <= 0;
          conv2d_4_col_select <= cparam_conv2d_4_col_select_initval;
          conv2d_4_filter_page_comp_offset_buf <= conv2d_4_filter_page_comp_offset;
          conv2d_4_act_page_comp_offset_buf_0 <= conv2d_4_act_page_comp_offset_0;
          conv2d_4_act_page_comp_offset_buf_1 <= conv2d_4_act_page_comp_offset_1;
          conv2d_4_act_page_comp_offset_buf_2 <= conv2d_4_act_page_comp_offset_2;
          conv2d_4_out_page_comp_offset_buf <= conv2d_4_out_page_comp_offset;
          conv2d_4_row_count_buf <= conv2d_4_row_count;
          conv2d_4_row_select_buf <= conv2d_4_row_select;
          conv2d_4_och_count_buf <= conv2d_4_och_count;
          conv2d_4_next_stream_num_ops <= (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)? cparam_conv2d_4_stream_num_ops_res : cparam_conv2d_4_stream_num_ops;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_2;
        end
        conv2d_4_comp_fsm_2: begin
          conv2d_4_stream_pad_masks <= { conv2d_4_stream_pad_mask_2_2, conv2d_4_stream_pad_mask_2_1, conv2d_4_stream_pad_mask_2_0, conv2d_4_stream_pad_mask_1_2, conv2d_4_stream_pad_mask_1_1, conv2d_4_stream_pad_mask_1_0, conv2d_4_stream_pad_mask_0_2, conv2d_4_stream_pad_mask_0_1, conv2d_4_stream_pad_mask_0_0 };
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_3;
        end
        conv2d_4_comp_fsm_3: begin
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          if(_stream_conv2d_4_stream_oready) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          end 
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
        end
        conv2d_4_comp_fsm_4: begin
          if(!_stream_conv2d_4_source_busy) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_5;
          end 
        end
        conv2d_4_comp_fsm_5: begin
          if(_stream_conv2d_4_busy) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_6;
          end 
        end
        conv2d_4_comp_fsm_6: begin
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_0 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_1 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_2 : 0)) begin
            conv2d_4_stream_act_local_0 <= conv2d_4_stream_act_local_0 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_0 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_1 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_2 : 0) begin
            conv2d_4_stream_act_local_0 <= conv2d_4_stream_act_local_0 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_0 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_0 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_0 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_3 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_4 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_5 : 0)) begin
            conv2d_4_stream_act_local_1 <= conv2d_4_stream_act_local_1 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_3 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_4 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_5 : 0) begin
            conv2d_4_stream_act_local_1 <= conv2d_4_stream_act_local_1 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_1 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_1 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_1 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_6 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_7 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_8 : 0)) begin
            conv2d_4_stream_act_local_2 <= conv2d_4_stream_act_local_2 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_6 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_7 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_8 : 0) begin
            conv2d_4_stream_act_local_2 <= conv2d_4_stream_act_local_2 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_2 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_2 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_2 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_9 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_10 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_11 : 0)) begin
            conv2d_4_stream_act_local_3 <= conv2d_4_stream_act_local_3 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_9 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_10 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_11 : 0) begin
            conv2d_4_stream_act_local_3 <= conv2d_4_stream_act_local_3 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_3 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_3 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_3 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_12 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_13 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_14 : 0)) begin
            conv2d_4_stream_act_local_4 <= conv2d_4_stream_act_local_4 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_12 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_13 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_14 : 0) begin
            conv2d_4_stream_act_local_4 <= conv2d_4_stream_act_local_4 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_4 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_4 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_4 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_15 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_16 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_17 : 0)) begin
            conv2d_4_stream_act_local_5 <= conv2d_4_stream_act_local_5 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_15 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_16 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_17 : 0) begin
            conv2d_4_stream_act_local_5 <= conv2d_4_stream_act_local_5 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_5 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_5 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_5 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_18 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_19 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_20 : 0)) begin
            conv2d_4_stream_act_local_6 <= conv2d_4_stream_act_local_6 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_18 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_19 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_20 : 0) begin
            conv2d_4_stream_act_local_6 <= conv2d_4_stream_act_local_6 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_6 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_6 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_6 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_21 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_22 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_23 : 0)) begin
            conv2d_4_stream_act_local_7 <= conv2d_4_stream_act_local_7 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_21 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_22 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_23 : 0) begin
            conv2d_4_stream_act_local_7 <= conv2d_4_stream_act_local_7 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_7 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_7 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_7 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_24 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_25 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_26 : 0)) begin
            conv2d_4_stream_act_local_8 <= conv2d_4_stream_act_local_8 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_24 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_25 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_26 : 0) begin
            conv2d_4_stream_act_local_8 <= conv2d_4_stream_act_local_8 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_8 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_8 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_8 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(cparam_conv2d_4_data_stationary == 0) begin
            conv2d_4_stream_out_local_col <= conv2d_4_stream_out_local_col + conv2d_4_next_stream_num_ops;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_col_count >= cparam_conv2d_4_max_col_count)) begin
            conv2d_4_stream_out_local_col <= 0;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            conv2d_4_stream_out_local_col <= conv2d_4_stream_out_local_col + cparam_conv2d_4_inc_out_laddr_col;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_col_count >= cparam_conv2d_4_max_col_count)) begin
            conv2d_4_stream_out_local_val <= conv2d_4_stream_out_local_val + conv2d_4_next_stream_num_ops;
            conv2d_4_stream_out_local_col <= 0;
          end 
          conv2d_4_col_count <= conv2d_4_col_count + cparam_conv2d_4_stride_col_par_col;
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_col_count <= 0;
          end 
          conv2d_4_col_select <= conv2d_4_col_select + cparam_conv2d_4_stride_col_mod_filter_num;
          if(conv2d_4_col_select + cparam_conv2d_4_stride_col_mod_filter_num >= 3) begin
            conv2d_4_col_select <= conv2d_4_col_select - cparam_conv2d_4_filter_num_col_minus_stride_col_mod;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_col_select <= cparam_conv2d_4_col_select_initval;
          end 
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_2;
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_336 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1)) begin
        _tmp_336 <= read_rtl_bank_335;
      end 
    end
  end

  localparam _stream_conv2d_4_source_7_source_pat_fsm_0_1 = 1;
  localparam _stream_conv2d_4_source_7_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_init;
    end else begin
      case(_stream_conv2d_4_source_7_source_pat_fsm_0)
        _stream_conv2d_4_source_7_source_pat_fsm_0_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_1;
          end 
        end
        _stream_conv2d_4_source_7_source_pat_fsm_0_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_init;
          end 
          if((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0) && (_source_stream_conv2d_4_source_7_pat_count_2 == 0) && (_source_stream_conv2d_4_source_7_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_2;
          end 
        end
        _stream_conv2d_4_source_7_source_pat_fsm_0_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_346 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2)) begin
        _tmp_346 <= read_rtl_bank_345;
      end 
    end
  end

  localparam _stream_conv2d_4_source_9_source_pat_fsm_1_1 = 1;
  localparam _stream_conv2d_4_source_9_source_pat_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_init;
    end else begin
      case(_stream_conv2d_4_source_9_source_pat_fsm_1)
        _stream_conv2d_4_source_9_source_pat_fsm_1_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_1;
          end 
        end
        _stream_conv2d_4_source_9_source_pat_fsm_1_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_init;
          end 
          if((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0) && (_source_stream_conv2d_4_source_9_pat_count_2 == 0) && (_source_stream_conv2d_4_source_9_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_2;
          end 
        end
        _stream_conv2d_4_source_9_source_pat_fsm_1_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_365 <= 0;
      _tmp_1366 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3)) begin
        _tmp_365 <= read_rtl_bank_364;
      end 
      if(_stream_matmul_23_stream_oready && _stream_matmul_23_source_7_source_ram_renable && (_stream_matmul_23_source_7_source_sel == 1)) begin
        _tmp_1366 <= read_rtl_bank_1365;
      end 
    end
  end

  localparam _stream_conv2d_4_source_20_source_pat_fsm_2_1 = 1;
  localparam _stream_conv2d_4_source_20_source_pat_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_init;
    end else begin
      case(_stream_conv2d_4_source_20_source_pat_fsm_2)
        _stream_conv2d_4_source_20_source_pat_fsm_2_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_1;
          end 
        end
        _stream_conv2d_4_source_20_source_pat_fsm_2_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_init;
          end 
          if((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0) && (_source_stream_conv2d_4_source_20_pat_count_2 == 0) && (_source_stream_conv2d_4_source_20_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_2;
          end 
        end
        _stream_conv2d_4_source_20_source_pat_fsm_2_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_374 <= 0;
      _tmp_1376 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4)) begin
        _tmp_374 <= read_rtl_bank_373;
      end 
      if(_stream_matmul_23_stream_oready && _stream_matmul_23_source_9_source_ram_renable && (_stream_matmul_23_source_9_source_sel == 2)) begin
        _tmp_1376 <= read_rtl_bank_1375;
      end 
    end
  end

  localparam _stream_conv2d_4_source_21_source_pat_fsm_3_1 = 1;
  localparam _stream_conv2d_4_source_21_source_pat_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_init;
    end else begin
      case(_stream_conv2d_4_source_21_source_pat_fsm_3)
        _stream_conv2d_4_source_21_source_pat_fsm_3_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_1;
          end 
        end
        _stream_conv2d_4_source_21_source_pat_fsm_3_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_init;
          end 
          if((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0) && (_source_stream_conv2d_4_source_21_pat_count_2 == 0) && (_source_stream_conv2d_4_source_21_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_2;
          end 
        end
        _stream_conv2d_4_source_21_source_pat_fsm_3_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_383 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5)) begin
        _tmp_383 <= read_rtl_bank_382;
      end 
    end
  end

  localparam _stream_conv2d_4_source_22_source_pat_fsm_4_1 = 1;
  localparam _stream_conv2d_4_source_22_source_pat_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_init;
    end else begin
      case(_stream_conv2d_4_source_22_source_pat_fsm_4)
        _stream_conv2d_4_source_22_source_pat_fsm_4_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_1;
          end 
        end
        _stream_conv2d_4_source_22_source_pat_fsm_4_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_init;
          end 
          if((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0) && (_source_stream_conv2d_4_source_22_pat_count_2 == 0) && (_source_stream_conv2d_4_source_22_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_2;
          end 
        end
        _stream_conv2d_4_source_22_source_pat_fsm_4_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_392 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6)) begin
        _tmp_392 <= read_rtl_bank_391;
      end 
    end
  end

  localparam _stream_conv2d_4_source_23_source_pat_fsm_5_1 = 1;
  localparam _stream_conv2d_4_source_23_source_pat_fsm_5_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_init;
    end else begin
      case(_stream_conv2d_4_source_23_source_pat_fsm_5)
        _stream_conv2d_4_source_23_source_pat_fsm_5_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_1;
          end 
        end
        _stream_conv2d_4_source_23_source_pat_fsm_5_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_init;
          end 
          if((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0) && (_source_stream_conv2d_4_source_23_pat_count_2 == 0) && (_source_stream_conv2d_4_source_23_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_2;
          end 
        end
        _stream_conv2d_4_source_23_source_pat_fsm_5_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_401 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7)) begin
        _tmp_401 <= read_rtl_bank_400;
      end 
    end
  end

  localparam _stream_conv2d_4_source_24_source_pat_fsm_6_1 = 1;
  localparam _stream_conv2d_4_source_24_source_pat_fsm_6_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_init;
    end else begin
      case(_stream_conv2d_4_source_24_source_pat_fsm_6)
        _stream_conv2d_4_source_24_source_pat_fsm_6_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_1;
          end 
        end
        _stream_conv2d_4_source_24_source_pat_fsm_6_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_init;
          end 
          if((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0) && (_source_stream_conv2d_4_source_24_pat_count_2 == 0) && (_source_stream_conv2d_4_source_24_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_2;
          end 
        end
        _stream_conv2d_4_source_24_source_pat_fsm_6_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_410 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8)) begin
        _tmp_410 <= read_rtl_bank_409;
      end 
    end
  end

  localparam _stream_conv2d_4_source_25_source_pat_fsm_7_1 = 1;
  localparam _stream_conv2d_4_source_25_source_pat_fsm_7_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_init;
    end else begin
      case(_stream_conv2d_4_source_25_source_pat_fsm_7)
        _stream_conv2d_4_source_25_source_pat_fsm_7_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_1;
          end 
        end
        _stream_conv2d_4_source_25_source_pat_fsm_7_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_init;
          end 
          if((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0) && (_source_stream_conv2d_4_source_25_pat_count_2 == 0) && (_source_stream_conv2d_4_source_25_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_2;
          end 
        end
        _stream_conv2d_4_source_25_source_pat_fsm_7_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_419 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9)) begin
        _tmp_419 <= read_rtl_bank_418;
      end 
    end
  end

  localparam _stream_conv2d_4_source_26_source_pat_fsm_8_1 = 1;
  localparam _stream_conv2d_4_source_26_source_pat_fsm_8_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_init;
    end else begin
      case(_stream_conv2d_4_source_26_source_pat_fsm_8)
        _stream_conv2d_4_source_26_source_pat_fsm_8_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_1;
          end 
        end
        _stream_conv2d_4_source_26_source_pat_fsm_8_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_init;
          end 
          if((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0) && (_source_stream_conv2d_4_source_26_pat_count_2 == 0) && (_source_stream_conv2d_4_source_26_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_2;
          end 
        end
        _stream_conv2d_4_source_26_source_pat_fsm_8_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_428 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10)) begin
        _tmp_428 <= read_rtl_bank_427;
      end 
    end
  end

  localparam _stream_conv2d_4_source_27_source_pat_fsm_9_1 = 1;
  localparam _stream_conv2d_4_source_27_source_pat_fsm_9_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_init;
    end else begin
      case(_stream_conv2d_4_source_27_source_pat_fsm_9)
        _stream_conv2d_4_source_27_source_pat_fsm_9_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_1;
          end 
        end
        _stream_conv2d_4_source_27_source_pat_fsm_9_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_init;
          end 
          if((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0) && (_source_stream_conv2d_4_source_27_pat_count_2 == 0) && (_source_stream_conv2d_4_source_27_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_2;
          end 
        end
        _stream_conv2d_4_source_27_source_pat_fsm_9_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_437 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11)) begin
        _tmp_437 <= read_rtl_bank_436;
      end 
    end
  end

  localparam _stream_conv2d_4_source_28_source_pat_fsm_10_1 = 1;
  localparam _stream_conv2d_4_source_28_source_pat_fsm_10_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_init;
    end else begin
      case(_stream_conv2d_4_source_28_source_pat_fsm_10)
        _stream_conv2d_4_source_28_source_pat_fsm_10_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_1;
          end 
        end
        _stream_conv2d_4_source_28_source_pat_fsm_10_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_init;
          end 
          if((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0) && (_source_stream_conv2d_4_source_28_pat_count_2 == 0) && (_source_stream_conv2d_4_source_28_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_2;
          end 
        end
        _stream_conv2d_4_source_28_source_pat_fsm_10_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_446 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12)) begin
        _tmp_446 <= read_rtl_bank_445;
      end 
    end
  end

  localparam _stream_conv2d_4_source_29_source_pat_fsm_11_1 = 1;
  localparam _stream_conv2d_4_source_29_source_pat_fsm_11_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_init;
    end else begin
      case(_stream_conv2d_4_source_29_source_pat_fsm_11)
        _stream_conv2d_4_source_29_source_pat_fsm_11_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_1;
          end 
        end
        _stream_conv2d_4_source_29_source_pat_fsm_11_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_init;
          end 
          if((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0) && (_source_stream_conv2d_4_source_29_pat_count_2 == 0) && (_source_stream_conv2d_4_source_29_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_2;
          end 
        end
        _stream_conv2d_4_source_29_source_pat_fsm_11_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_455 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13)) begin
        _tmp_455 <= read_rtl_bank_454;
      end 
    end
  end

  localparam _stream_conv2d_4_source_30_source_pat_fsm_12_1 = 1;
  localparam _stream_conv2d_4_source_30_source_pat_fsm_12_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_init;
    end else begin
      case(_stream_conv2d_4_source_30_source_pat_fsm_12)
        _stream_conv2d_4_source_30_source_pat_fsm_12_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_1;
          end 
        end
        _stream_conv2d_4_source_30_source_pat_fsm_12_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_init;
          end 
          if((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0) && (_source_stream_conv2d_4_source_30_pat_count_2 == 0) && (_source_stream_conv2d_4_source_30_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_2;
          end 
        end
        _stream_conv2d_4_source_30_source_pat_fsm_12_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_464 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14)) begin
        _tmp_464 <= read_rtl_bank_463;
      end 
    end
  end

  localparam _stream_conv2d_4_source_31_source_pat_fsm_13_1 = 1;
  localparam _stream_conv2d_4_source_31_source_pat_fsm_13_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_init;
    end else begin
      case(_stream_conv2d_4_source_31_source_pat_fsm_13)
        _stream_conv2d_4_source_31_source_pat_fsm_13_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_1;
          end 
        end
        _stream_conv2d_4_source_31_source_pat_fsm_13_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_init;
          end 
          if((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0) && (_source_stream_conv2d_4_source_31_pat_count_2 == 0) && (_source_stream_conv2d_4_source_31_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_2;
          end 
        end
        _stream_conv2d_4_source_31_source_pat_fsm_13_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_473 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15)) begin
        _tmp_473 <= read_rtl_bank_472;
      end 
    end
  end

  localparam _stream_conv2d_4_source_32_source_pat_fsm_14_1 = 1;
  localparam _stream_conv2d_4_source_32_source_pat_fsm_14_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_init;
    end else begin
      case(_stream_conv2d_4_source_32_source_pat_fsm_14)
        _stream_conv2d_4_source_32_source_pat_fsm_14_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_1;
          end 
        end
        _stream_conv2d_4_source_32_source_pat_fsm_14_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_init;
          end 
          if((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0) && (_source_stream_conv2d_4_source_32_pat_count_2 == 0) && (_source_stream_conv2d_4_source_32_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_2;
          end 
        end
        _stream_conv2d_4_source_32_source_pat_fsm_14_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_482 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16)) begin
        _tmp_482 <= read_rtl_bank_481;
      end 
    end
  end

  localparam _stream_conv2d_4_source_33_source_pat_fsm_15_1 = 1;
  localparam _stream_conv2d_4_source_33_source_pat_fsm_15_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_init;
    end else begin
      case(_stream_conv2d_4_source_33_source_pat_fsm_15)
        _stream_conv2d_4_source_33_source_pat_fsm_15_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_1;
          end 
        end
        _stream_conv2d_4_source_33_source_pat_fsm_15_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_init;
          end 
          if((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0) && (_source_stream_conv2d_4_source_33_pat_count_2 == 0) && (_source_stream_conv2d_4_source_33_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_2;
          end 
        end
        _stream_conv2d_4_source_33_source_pat_fsm_15_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_491 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17)) begin
        _tmp_491 <= read_rtl_bank_490;
      end 
    end
  end

  localparam _stream_conv2d_4_source_34_source_pat_fsm_16_1 = 1;
  localparam _stream_conv2d_4_source_34_source_pat_fsm_16_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_init;
    end else begin
      case(_stream_conv2d_4_source_34_source_pat_fsm_16)
        _stream_conv2d_4_source_34_source_pat_fsm_16_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_1;
          end 
        end
        _stream_conv2d_4_source_34_source_pat_fsm_16_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_init;
          end 
          if((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0) && (_source_stream_conv2d_4_source_34_pat_count_2 == 0) && (_source_stream_conv2d_4_source_34_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_2;
          end 
        end
        _stream_conv2d_4_source_34_source_pat_fsm_16_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_500 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18)) begin
        _tmp_500 <= read_rtl_bank_499;
      end 
    end
  end

  localparam _stream_conv2d_4_source_35_source_pat_fsm_17_1 = 1;
  localparam _stream_conv2d_4_source_35_source_pat_fsm_17_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_init;
    end else begin
      case(_stream_conv2d_4_source_35_source_pat_fsm_17)
        _stream_conv2d_4_source_35_source_pat_fsm_17_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_1;
          end 
        end
        _stream_conv2d_4_source_35_source_pat_fsm_17_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_init;
          end 
          if((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0) && (_source_stream_conv2d_4_source_35_pat_count_2 == 0) && (_source_stream_conv2d_4_source_35_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_2;
          end 
        end
        _stream_conv2d_4_source_35_source_pat_fsm_17_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_509 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19)) begin
        _tmp_509 <= read_rtl_bank_508;
      end 
    end
  end

  localparam _stream_conv2d_4_source_36_source_pat_fsm_18_1 = 1;
  localparam _stream_conv2d_4_source_36_source_pat_fsm_18_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_init;
    end else begin
      case(_stream_conv2d_4_source_36_source_pat_fsm_18)
        _stream_conv2d_4_source_36_source_pat_fsm_18_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_1;
          end 
        end
        _stream_conv2d_4_source_36_source_pat_fsm_18_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_init;
          end 
          if((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0) && (_source_stream_conv2d_4_source_36_pat_count_2 == 0) && (_source_stream_conv2d_4_source_36_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_2;
          end 
        end
        _stream_conv2d_4_source_36_source_pat_fsm_18_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_518 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20)) begin
        _tmp_518 <= read_rtl_bank_517;
      end 
    end
  end

  localparam _stream_conv2d_4_source_37_source_pat_fsm_19_1 = 1;
  localparam _stream_conv2d_4_source_37_source_pat_fsm_19_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_init;
    end else begin
      case(_stream_conv2d_4_source_37_source_pat_fsm_19)
        _stream_conv2d_4_source_37_source_pat_fsm_19_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_1;
          end 
        end
        _stream_conv2d_4_source_37_source_pat_fsm_19_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_init;
          end 
          if((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0) && (_source_stream_conv2d_4_source_37_pat_count_2 == 0) && (_source_stream_conv2d_4_source_37_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_2;
          end 
        end
        _stream_conv2d_4_source_37_source_pat_fsm_19_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_sink_50_sink_fsm_20_1 = 1;
  localparam _stream_conv2d_4_sink_50_sink_fsm_20_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_sink_50_sink_fsm_20 <= _stream_conv2d_4_sink_50_sink_fsm_20_init;
    end else begin
      case(_stream_conv2d_4_sink_50_sink_fsm_20)
        _stream_conv2d_4_sink_50_sink_fsm_20_init: begin
          if(_stream_conv2d_4_sink_start && _stream_conv2d_4_sink_50_sink_mode & 5'b1 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_sink_50_sink_fsm_20 <= _stream_conv2d_4_sink_50_sink_fsm_20_1;
          end 
        end
        _stream_conv2d_4_sink_50_sink_fsm_20_1: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_sink_50_sink_fsm_20 <= _stream_conv2d_4_sink_50_sink_fsm_20_2;
          end 
        end
        _stream_conv2d_4_sink_50_sink_fsm_20_2: begin
          if(stream_conv2d_4_sink_51_data && (_stream_conv2d_4_sink_50_sink_count == 1) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_sink_50_sink_fsm_20 <= _stream_conv2d_4_sink_50_sink_fsm_20_init;
          end 
          if(_stream_conv2d_4_sink_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_sink_50_sink_fsm_20 <= _stream_conv2d_4_sink_50_sink_fsm_20_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_write_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_write_req_fsm <= _maxi_write_req_fsm_init;
      _maxi_write_cont <= 0;
    end else begin
      case(_maxi_write_req_fsm)
        _maxi_write_req_fsm_init: begin
          if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full) begin
            _maxi_write_req_fsm <= _maxi_write_req_fsm_1;
          end 
        end
        _maxi_write_req_fsm_1: begin
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) begin
            _maxi_write_cont <= 1;
          end 
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6) && (_maxi_write_global_size == 0)) begin
            _maxi_write_cont <= 0;
          end 
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) begin
            _maxi_write_req_fsm <= _maxi_write_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_write_data_fsm_1 = 1;
  localparam _maxi_write_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
    end else begin
      case(_maxi_write_data_fsm)
        _maxi_write_data_fsm_init: begin
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
        end
        _maxi_write_data_fsm_1: begin
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
        end
        _maxi_write_data_fsm_2: begin
          if((_maxi_write_op_sel_buf == 1) && read_burst_packed_rvalid_1169 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_packed_rlast_1170) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
          if((_maxi_write_op_sel_buf == 2) && read_burst_rvalid_1301 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_rlast_1302) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
          if((_maxi_write_op_sel_buf == 3) && read_burst_rvalid_2012 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_rlast_2013) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_packed_fsm_24_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_packed_fsm_24 <= read_burst_packed_fsm_24_init;
      read_burst_packed_addr_1166 <= 0;
      read_burst_packed_stride_1167 <= 0;
      read_burst_packed_length_1168 <= 0;
      read_burst_packed_rvalid_1169 <= 0;
      read_burst_packed_rlast_1170 <= 0;
    end else begin
      case(read_burst_packed_fsm_24)
        read_burst_packed_fsm_24_init: begin
          read_burst_packed_addr_1166 <= _maxi_write_local_addr_buf;
          read_burst_packed_stride_1167 <= _maxi_write_local_stride_buf;
          read_burst_packed_length_1168 <= _maxi_write_size_buf;
          read_burst_packed_rvalid_1169 <= 0;
          read_burst_packed_rlast_1170 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 1) && (_maxi_write_size_buf > 0)) begin
            read_burst_packed_fsm_24 <= read_burst_packed_fsm_24_1;
          end 
        end
        read_burst_packed_fsm_24_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1168 > 0)) begin
            read_burst_packed_addr_1166 <= read_burst_packed_addr_1166 + read_burst_packed_stride_1167;
            read_burst_packed_length_1168 <= read_burst_packed_length_1168 - 1;
            read_burst_packed_rvalid_1169 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1168 <= 1)) begin
            read_burst_packed_rlast_1170 <= 1;
          end 
          if(read_burst_packed_rlast_1170 && read_burst_packed_rvalid_1169 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_rvalid_1169 <= 0;
            read_burst_packed_rlast_1170 <= 0;
          end 
          if(0) begin
            read_burst_packed_rvalid_1169 <= 0;
            read_burst_packed_rlast_1170 <= 0;
          end 
          if(read_burst_packed_rlast_1170 && read_burst_packed_rvalid_1169 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_fsm_24 <= read_burst_packed_fsm_24_init;
          end 
          if(0) begin
            read_burst_packed_fsm_24 <= read_burst_packed_fsm_24_init;
          end 
        end
      endcase
    end
  end

  localparam control_max_pool_serial_6_1 = 1;
  localparam control_max_pool_serial_6_2 = 2;
  localparam control_max_pool_serial_6_3 = 3;
  localparam control_max_pool_serial_6_4 = 4;
  localparam control_max_pool_serial_6_5 = 5;
  localparam control_max_pool_serial_6_6 = 6;
  localparam control_max_pool_serial_6_7 = 7;
  localparam control_max_pool_serial_6_8 = 8;
  localparam control_max_pool_serial_6_9 = 9;
  localparam control_max_pool_serial_6_10 = 10;
  localparam control_max_pool_serial_6_11 = 11;
  localparam control_max_pool_serial_6_12 = 12;
  localparam control_max_pool_serial_6_13 = 13;
  localparam control_max_pool_serial_6_14 = 14;
  localparam control_max_pool_serial_6_15 = 15;
  localparam control_max_pool_serial_6_16 = 16;
  localparam control_max_pool_serial_6_17 = 17;
  localparam control_max_pool_serial_6_18 = 18;
  localparam control_max_pool_serial_6_19 = 19;

  always @(posedge CLK) begin
    if(RST) begin
      control_max_pool_serial_6 <= control_max_pool_serial_6_init;
      _control_max_pool_serial_6_called <= 0;
      max_pool_serial_6_act_base_offset_row <= 0;
      max_pool_serial_6_act_base_offset_bat <= 0;
      max_pool_serial_6_act_page <= 0;
      max_pool_serial_6_act_page_comp_offset <= 0;
      max_pool_serial_6_act_page_dma_offset <= 0;
      max_pool_serial_6_out_base_offset_row <= 0;
      max_pool_serial_6_out_base_offset_bat <= 0;
      max_pool_serial_6_out_page <= 0;
      max_pool_serial_6_out_page_comp_offset <= 0;
      max_pool_serial_6_out_page_dma_offset <= 0;
      max_pool_serial_6_row_count <= 0;
      max_pool_serial_6_bat_count <= 0;
      max_pool_serial_6_prev_row_count <= 0;
      max_pool_serial_6_prev_bat_count <= 0;
      max_pool_serial_6_skip_read_act <= 0;
      max_pool_serial_6_skip_comp <= 0;
      max_pool_serial_6_skip_write_out <= 0;
      max_pool_serial_6_out_count <= 0;
    end else begin
      case(control_max_pool_serial_6)
        control_max_pool_serial_6_init: begin
          if(main_fsm == 18) begin
            _control_max_pool_serial_6_called <= 1;
          end 
          if(main_fsm == 35) begin
            _control_max_pool_serial_6_called <= 1;
          end 
          if(main_fsm == 52) begin
            _control_max_pool_serial_6_called <= 1;
          end 
          if(main_fsm == 18) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_1;
          end 
          if(main_fsm == 35) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_1;
          end 
          if(main_fsm == 52) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_1;
          end 
        end
        control_max_pool_serial_6_1: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_2;
        end
        control_max_pool_serial_6_2: begin
          max_pool_serial_6_act_base_offset_row <= 0;
          max_pool_serial_6_act_base_offset_bat <= 0;
          max_pool_serial_6_act_page <= 0;
          max_pool_serial_6_act_page_comp_offset <= 0;
          max_pool_serial_6_act_page_dma_offset <= 0;
          max_pool_serial_6_out_base_offset_row <= 0;
          max_pool_serial_6_out_base_offset_bat <= 0;
          max_pool_serial_6_out_page <= 0;
          max_pool_serial_6_out_page_comp_offset <= 0;
          max_pool_serial_6_out_page_dma_offset <= 0;
          max_pool_serial_6_row_count <= 0;
          max_pool_serial_6_bat_count <= 0;
          max_pool_serial_6_prev_row_count <= 0;
          max_pool_serial_6_prev_bat_count <= 0;
          max_pool_serial_6_skip_read_act <= 0;
          max_pool_serial_6_skip_comp <= 0;
          max_pool_serial_6_skip_write_out <= 1;
          max_pool_serial_6_out_count <= 0;
          control_max_pool_serial_6 <= control_max_pool_serial_6_3;
        end
        control_max_pool_serial_6_3: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_4;
          if(max_pool_serial_6_skip_read_act) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_11;
          end 
        end
        control_max_pool_serial_6_4: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_5;
          if(max_pool_serial_6_dma_pad_mask_0) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_7;
          end 
        end
        control_max_pool_serial_6_5: begin
          if(_maxi_read_req_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_6;
          end 
        end
        control_max_pool_serial_6_6: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_7;
          end 
        end
        control_max_pool_serial_6_7: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_8;
          if(max_pool_serial_6_dma_pad_mask_1) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_10;
          end 
        end
        control_max_pool_serial_6_8: begin
          if(_maxi_read_req_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_9;
          end 
        end
        control_max_pool_serial_6_9: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_10;
          end 
        end
        control_max_pool_serial_6_10: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_11;
        end
        control_max_pool_serial_6_11: begin
          if(_maxi_write_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_12;
          end 
        end
        control_max_pool_serial_6_12: begin
          if(max_pool_serial_6_comp_fsm == 0) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_13;
          end 
        end
        control_max_pool_serial_6_13: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_14;
          if(max_pool_serial_6_skip_write_out) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_17;
          end 
        end
        control_max_pool_serial_6_14: begin
          if(max_pool_serial_6_comp_count >= max_pool_serial_6_out_count + cparam_max_pool_serial_6_out_write_size) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_15;
          end 
        end
        control_max_pool_serial_6_15: begin
          if(_maxi_write_req_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_16;
          end 
        end
        control_max_pool_serial_6_16: begin
          max_pool_serial_6_out_count <= max_pool_serial_6_out_count + cparam_max_pool_serial_6_out_write_size;
          control_max_pool_serial_6 <= control_max_pool_serial_6_17;
        end
        control_max_pool_serial_6_17: begin
          max_pool_serial_6_act_base_offset_row <= max_pool_serial_6_act_base_offset_row + cparam_max_pool_serial_6_act_row_step;
          if(max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) begin
            max_pool_serial_6_act_base_offset_row <= 0;
            max_pool_serial_6_act_base_offset_bat <= max_pool_serial_6_act_base_offset_bat + cparam_max_pool_serial_6_act_bat_step;
          end 
          if((max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_act_base_offset_bat <= 0;
          end 
          max_pool_serial_6_row_count <= max_pool_serial_6_row_count + cparam_max_pool_serial_6_stride_row;
          if(max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) begin
            max_pool_serial_6_row_count <= 0;
            max_pool_serial_6_bat_count <= max_pool_serial_6_bat_count + 1;
          end 
          if((max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_bat_count <= 0;
          end 
          if(!max_pool_serial_6_act_page) begin
            max_pool_serial_6_act_page_comp_offset <= 2048;
            max_pool_serial_6_act_page_dma_offset <= 2048;
            max_pool_serial_6_act_page <= 1;
          end 
          if(max_pool_serial_6_act_page) begin
            max_pool_serial_6_act_page_comp_offset <= 0;
            max_pool_serial_6_act_page_dma_offset <= 0;
            max_pool_serial_6_act_page <= 0;
          end 
          if(!max_pool_serial_6_skip_write_out) begin
            max_pool_serial_6_out_base_offset_row <= max_pool_serial_6_out_base_offset_row + cparam_max_pool_serial_6_out_row_step;
          end 
          if(!max_pool_serial_6_skip_write_out && (max_pool_serial_6_prev_row_count >= cparam_max_pool_serial_6_max_row_count)) begin
            max_pool_serial_6_out_base_offset_row <= 0;
            max_pool_serial_6_out_base_offset_bat <= max_pool_serial_6_out_base_offset_bat + cparam_max_pool_serial_6_out_bat_step;
          end 
          if(!max_pool_serial_6_skip_write_out && (max_pool_serial_6_prev_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_prev_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_out_base_offset_bat <= 0;
          end 
          if(!max_pool_serial_6_out_page) begin
            max_pool_serial_6_out_page_comp_offset <= 512;
            max_pool_serial_6_out_page_dma_offset <= 0;
            max_pool_serial_6_out_page <= 1;
          end 
          if(max_pool_serial_6_out_page) begin
            max_pool_serial_6_out_page_comp_offset <= 0;
            max_pool_serial_6_out_page_dma_offset <= 512;
            max_pool_serial_6_out_page <= 0;
          end 
          max_pool_serial_6_prev_row_count <= max_pool_serial_6_row_count;
          max_pool_serial_6_prev_bat_count <= max_pool_serial_6_bat_count;
          if((max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_skip_read_act <= 1;
          end 
          if((max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_skip_comp <= 1;
          end 
          if(max_pool_serial_6_skip_write_out && (max_pool_serial_6_prev_row_count == 0) && (max_pool_serial_6_prev_bat_count == 0)) begin
            max_pool_serial_6_skip_write_out <= 0;
          end 
          control_max_pool_serial_6 <= control_max_pool_serial_6_3;
          if(!max_pool_serial_6_skip_write_out && (max_pool_serial_6_prev_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_prev_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_18;
          end 
        end
        control_max_pool_serial_6_18: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_19;
          end 
        end
        control_max_pool_serial_6_19: begin
          if(main_fsm == 21) begin
            _control_max_pool_serial_6_called <= 0;
          end 
          if(main_fsm == 38) begin
            _control_max_pool_serial_6_called <= 0;
          end 
          if(main_fsm == 55) begin
            _control_max_pool_serial_6_called <= 0;
          end 
          if(main_fsm == 21) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_init;
          end 
          if(main_fsm == 38) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_init;
          end 
          if(main_fsm == 55) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_25_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_25 <= write_burst_fsm_25_init;
      write_burst_addr_1182 <= 0;
      write_burst_stride_1183 <= 0;
      write_burst_length_1184 <= 0;
      write_burst_done_1185 <= 0;
    end else begin
      case(write_burst_fsm_25)
        write_burst_fsm_25_init: begin
          write_burst_addr_1182 <= _maxi_read_local_addr_buf;
          write_burst_stride_1183 <= _maxi_read_local_stride_buf;
          write_burst_length_1184 <= _maxi_read_local_size_buf;
          write_burst_done_1185 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 7) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_25 <= write_burst_fsm_25_1;
          end 
        end
        write_burst_fsm_25_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_1182 <= write_burst_addr_1182 + write_burst_stride_1183;
            write_burst_length_1184 <= write_burst_length_1184 - 1;
            write_burst_done_1185 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_1184 <= 1)) begin
            write_burst_done_1185 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_1185 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_1184 <= 1)) begin
            write_burst_fsm_25 <= write_burst_fsm_25_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_25 <= write_burst_fsm_25_init;
          end 
          if(0) begin
            write_burst_fsm_25 <= write_burst_fsm_25_init;
          end 
        end
      endcase
    end
  end

  localparam max_pool_serial_6_comp_fsm_1 = 1;
  localparam max_pool_serial_6_comp_fsm_2 = 2;
  localparam max_pool_serial_6_comp_fsm_3 = 3;
  localparam max_pool_serial_6_comp_fsm_4 = 4;
  localparam max_pool_serial_6_comp_fsm_5 = 5;
  localparam max_pool_serial_6_comp_fsm_6 = 6;
  localparam max_pool_serial_6_comp_fsm_7 = 7;

  always @(posedge CLK) begin
    if(RST) begin
      max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_init;
      max_pool_serial_6_stream_act_local <= 0;
      max_pool_serial_6_stream_out_local <= 0;
      max_pool_serial_6_col_count <= 0;
      max_pool_serial_6_act_page_comp_offset_buf <= 0;
      max_pool_serial_6_out_page_comp_offset_buf <= 0;
      max_pool_serial_6_row_count_buf <= 0;
      max_pool_serial_6_stream_pad_masks <= 0;
      max_pool_serial_6_comp_count <= 0;
    end else begin
      if(control_max_pool_serial_6 == 2) begin
        max_pool_serial_6_comp_count <= 0;
      end 
      if(_stream_max_pool_serial_6_sink_stop) begin
        max_pool_serial_6_comp_count <= max_pool_serial_6_comp_count + cparam_max_pool_serial_6_inc_out_laddr;
      end 
      case(max_pool_serial_6_comp_fsm)
        max_pool_serial_6_comp_fsm_init: begin
          if((control_max_pool_serial_6 == 12) && !max_pool_serial_6_skip_comp) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_1;
          end 
        end
        max_pool_serial_6_comp_fsm_1: begin
          max_pool_serial_6_stream_act_local <= cparam_max_pool_serial_6_local_pad_offset;
          max_pool_serial_6_stream_out_local <= 0;
          max_pool_serial_6_col_count <= 0;
          max_pool_serial_6_act_page_comp_offset_buf <= max_pool_serial_6_act_page_comp_offset;
          max_pool_serial_6_out_page_comp_offset_buf <= max_pool_serial_6_out_page_comp_offset;
          max_pool_serial_6_row_count_buf <= max_pool_serial_6_row_count;
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_2;
        end
        max_pool_serial_6_comp_fsm_2: begin
          max_pool_serial_6_stream_pad_masks <= { max_pool_serial_6_stream_pad_mask_1_1, max_pool_serial_6_stream_pad_mask_1_0, max_pool_serial_6_stream_pad_mask_0_1, max_pool_serial_6_stream_pad_mask_0_0 };
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_3;
        end
        max_pool_serial_6_comp_fsm_3: begin
          if(!_stream_max_pool_serial_6_source_busy) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_4;
          end 
        end
        max_pool_serial_6_comp_fsm_4: begin
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_5;
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_5;
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_5;
          if(_stream_max_pool_serial_6_stream_oready) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_5;
          end 
        end
        max_pool_serial_6_comp_fsm_5: begin
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_6;
        end
        max_pool_serial_6_comp_fsm_6: begin
          if(_stream_max_pool_serial_6_busy) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_7;
          end 
        end
        max_pool_serial_6_comp_fsm_7: begin
          max_pool_serial_6_stream_act_local <= max_pool_serial_6_stream_act_local + cparam_max_pool_serial_6_inc_act_laddr;
          if(max_pool_serial_6_col_count >= cparam_max_pool_serial_6_max_col_count) begin
            max_pool_serial_6_stream_act_local <= cparam_max_pool_serial_6_local_pad_offset;
          end 
          max_pool_serial_6_stream_out_local <= max_pool_serial_6_stream_out_local + cparam_max_pool_serial_6_inc_out_laddr;
          if(max_pool_serial_6_col_count >= cparam_max_pool_serial_6_max_col_count) begin
            max_pool_serial_6_stream_out_local <= 0;
          end 
          max_pool_serial_6_col_count <= max_pool_serial_6_col_count + cparam_max_pool_serial_6_stride_col;
          if(max_pool_serial_6_col_count >= cparam_max_pool_serial_6_max_col_count) begin
            max_pool_serial_6_col_count <= 0;
          end 
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_2;
          if(max_pool_serial_6_col_count >= cparam_max_pool_serial_6_max_col_count) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_serial_6_source_1_source_pat_fsm_0_1 = 1;
  localparam _stream_max_pool_serial_6_source_1_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init;
    end else begin
      case(_stream_max_pool_serial_6_source_1_source_pat_fsm_0)
        _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init: begin
          if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_1;
          end 
        end
        _stream_max_pool_serial_6_source_1_source_pat_fsm_0_1: begin
          if(_stream_max_pool_serial_6_source_stop && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init;
          end 
          if((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_2 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_3 == 0) && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_2;
          end 
        end
        _stream_max_pool_serial_6_source_1_source_pat_fsm_0_2: begin
          if(_stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_serial_6_sink_6_sink_fsm_1_1 = 1;
  localparam _stream_max_pool_serial_6_sink_6_sink_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_6_sink_6_sink_fsm_1 <= _stream_max_pool_serial_6_sink_6_sink_fsm_1_init;
    end else begin
      case(_stream_max_pool_serial_6_sink_6_sink_fsm_1)
        _stream_max_pool_serial_6_sink_6_sink_fsm_1_init: begin
          if(_stream_max_pool_serial_6_sink_start && _stream_max_pool_serial_6_sink_6_sink_mode & 5'b1 && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_sink_6_sink_fsm_1 <= _stream_max_pool_serial_6_sink_6_sink_fsm_1_1;
          end 
        end
        _stream_max_pool_serial_6_sink_6_sink_fsm_1_1: begin
          if(_stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_sink_6_sink_fsm_1 <= _stream_max_pool_serial_6_sink_6_sink_fsm_1_2;
          end 
        end
        _stream_max_pool_serial_6_sink_6_sink_fsm_1_2: begin
          if(stream_max_pool_serial_6_sink_7_data && (_stream_max_pool_serial_6_sink_6_sink_count == 1) && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_sink_6_sink_fsm_1 <= _stream_max_pool_serial_6_sink_6_sink_fsm_1_init;
          end 
          if(_stream_max_pool_serial_6_sink_stop && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_sink_6_sink_fsm_1 <= _stream_max_pool_serial_6_sink_6_sink_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_fsm_26_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_fsm_26 <= read_burst_fsm_26_init;
      read_burst_addr_1298 <= 0;
      read_burst_stride_1299 <= 0;
      read_burst_length_1300 <= 0;
      read_burst_rvalid_1301 <= 0;
      read_burst_rlast_1302 <= 0;
    end else begin
      case(read_burst_fsm_26)
        read_burst_fsm_26_init: begin
          read_burst_addr_1298 <= _maxi_write_local_addr_buf;
          read_burst_stride_1299 <= _maxi_write_local_stride_buf;
          read_burst_length_1300 <= _maxi_write_size_buf;
          read_burst_rvalid_1301 <= 0;
          read_burst_rlast_1302 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 2) && (_maxi_write_size_buf > 0)) begin
            read_burst_fsm_26 <= read_burst_fsm_26_1;
          end 
        end
        read_burst_fsm_26_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_1300 > 0)) begin
            read_burst_addr_1298 <= read_burst_addr_1298 + read_burst_stride_1299;
            read_burst_length_1300 <= read_burst_length_1300 - 1;
            read_burst_rvalid_1301 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_1300 <= 1)) begin
            read_burst_rlast_1302 <= 1;
          end 
          if(read_burst_rlast_1302 && read_burst_rvalid_1301 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_rvalid_1301 <= 0;
            read_burst_rlast_1302 <= 0;
          end 
          if(0) begin
            read_burst_rvalid_1301 <= 0;
            read_burst_rlast_1302 <= 0;
          end 
          if(read_burst_rlast_1302 && read_burst_rvalid_1301 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_fsm_26 <= read_burst_fsm_26_init;
          end 
          if(0) begin
            read_burst_fsm_26 <= read_burst_fsm_26_init;
          end 
        end
      endcase
    end
  end

  localparam control_matmul_23_1 = 1;
  localparam control_matmul_23_2 = 2;
  localparam control_matmul_23_3 = 3;
  localparam control_matmul_23_4 = 4;
  localparam control_matmul_23_5 = 5;
  localparam control_matmul_23_6 = 6;
  localparam control_matmul_23_7 = 7;
  localparam control_matmul_23_8 = 8;
  localparam control_matmul_23_9 = 9;
  localparam control_matmul_23_10 = 10;
  localparam control_matmul_23_11 = 11;
  localparam control_matmul_23_12 = 12;
  localparam control_matmul_23_13 = 13;
  localparam control_matmul_23_14 = 14;
  localparam control_matmul_23_15 = 15;
  localparam control_matmul_23_16 = 16;
  localparam control_matmul_23_17 = 17;
  localparam control_matmul_23_18 = 18;
  localparam control_matmul_23_19 = 19;
  localparam control_matmul_23_20 = 20;
  localparam control_matmul_23_21 = 21;
  localparam control_matmul_23_22 = 22;
  localparam control_matmul_23_23 = 23;
  localparam control_matmul_23_24 = 24;
  localparam control_matmul_23_25 = 25;
  localparam control_matmul_23_26 = 26;
  localparam control_matmul_23_27 = 27;
  localparam control_matmul_23_28 = 28;

  always @(posedge CLK) begin
    if(RST) begin
      control_matmul_23 <= control_matmul_23_init;
      _control_matmul_23_called <= 0;
      matmul_23_filter_base_offset <= 0;
      matmul_23_filter_page_comp_offset <= 0;
      matmul_23_filter_page_dma_offset <= 0;
      matmul_23_act_base_offset_row <= 0;
      matmul_23_act_base_offset_bat <= 0;
      matmul_23_dma_flag_0 <= 0;
      matmul_23_act_page_comp_offset_0 <= 0;
      matmul_23_act_page_dma_offset_0 <= 0;
      matmul_23_out_base_offset_val <= 0;
      matmul_23_out_base_offset_col <= 0;
      matmul_23_out_base_offset_row <= 0;
      matmul_23_out_base_offset_bat <= 0;
      matmul_23_out_base_offset_och <= 0;
      matmul_23_out_page <= 0;
      matmul_23_out_page_comp_offset <= 0;
      matmul_23_out_page_dma_offset <= 0;
      matmul_23_out_laddr_offset <= 0;
      matmul_23_sync_out_count <= 0;
      matmul_23_write_count <= 0;
      matmul_23_next_out_write_size <= 0;
      matmul_23_row_count <= 0;
      matmul_23_bat_count <= 0;
      matmul_23_och_count <= 0;
      matmul_23_row_select <= 0;
      matmul_23_prev_row_count <= 0;
      matmul_23_prev_bat_count <= 0;
      matmul_23_prev_och_count <= 0;
      matmul_23_prev_row_select <= 0;
      matmul_23_out_col_count <= 0;
      matmul_23_out_row_count <= 0;
      matmul_23_out_ram_select <= 0;
      matmul_23_skip_read_filter <= 0;
      matmul_23_skip_read_act <= 0;
      matmul_23_skip_comp <= 0;
      matmul_23_skip_write_out <= 1;
    end else begin
      case(control_matmul_23)
        control_matmul_23_init: begin
          if(main_fsm == 64) begin
            _control_matmul_23_called <= 1;
          end 
          if(main_fsm == 74) begin
            _control_matmul_23_called <= 1;
          end 
          if(main_fsm == 64) begin
            control_matmul_23 <= control_matmul_23_1;
          end 
          if(main_fsm == 74) begin
            control_matmul_23 <= control_matmul_23_1;
          end 
        end
        control_matmul_23_1: begin
          control_matmul_23 <= control_matmul_23_2;
        end
        control_matmul_23_2: begin
          matmul_23_filter_base_offset <= 0;
          matmul_23_filter_page_comp_offset <= 0;
          matmul_23_filter_page_dma_offset <= 0;
          matmul_23_act_base_offset_row <= 0;
          matmul_23_act_base_offset_bat <= 0;
          matmul_23_dma_flag_0 <= 1;
          matmul_23_act_page_comp_offset_0 <= 0;
          matmul_23_act_page_dma_offset_0 <= 0;
          matmul_23_out_base_offset_val <= 0;
          matmul_23_out_base_offset_col <= 0;
          matmul_23_out_base_offset_row <= 0;
          matmul_23_out_base_offset_bat <= 0;
          matmul_23_out_base_offset_och <= 0;
          matmul_23_out_page <= 0;
          matmul_23_out_page_comp_offset <= 0;
          matmul_23_out_page_dma_offset <= 0;
          matmul_23_out_laddr_offset <= 0;
          matmul_23_sync_out_count <= 0;
          matmul_23_write_count <= 0;
          matmul_23_next_out_write_size <= (cparam_matmul_23_max_och_count == 0)? cparam_matmul_23_out_write_size_res : cparam_matmul_23_out_write_size;
          matmul_23_row_count <= 0;
          matmul_23_bat_count <= 0;
          matmul_23_och_count <= 0;
          matmul_23_row_select <= 0;
          matmul_23_prev_row_count <= 0;
          matmul_23_prev_bat_count <= 0;
          matmul_23_prev_och_count <= 0;
          matmul_23_prev_row_select <= 0;
          matmul_23_out_col_count <= 0;
          matmul_23_out_row_count <= 0;
          matmul_23_out_ram_select <= 0;
          matmul_23_skip_read_filter <= 0;
          matmul_23_skip_read_act <= 0;
          matmul_23_skip_comp <= 0;
          matmul_23_skip_write_out <= 1;
          if(_maxi_read_req_idle) begin
            control_matmul_23 <= control_matmul_23_3;
          end 
        end
        control_matmul_23_3: begin
          if(_maxi_read_idle) begin
            control_matmul_23 <= control_matmul_23_4;
          end 
        end
        control_matmul_23_4: begin
          if(_maxi_read_req_idle) begin
            control_matmul_23 <= control_matmul_23_5;
          end 
        end
        control_matmul_23_5: begin
          if(_maxi_read_idle) begin
            control_matmul_23 <= control_matmul_23_6;
          end 
        end
        control_matmul_23_6: begin
          if(cparam_matmul_23_data_stationary == 0) begin
            control_matmul_23 <= control_matmul_23_7;
          end 
          if(cparam_matmul_23_data_stationary == 1) begin
            control_matmul_23 <= control_matmul_23_12;
          end 
        end
        control_matmul_23_7: begin
          control_matmul_23 <= control_matmul_23_8;
          if(matmul_23_skip_read_filter) begin
            control_matmul_23 <= control_matmul_23_11;
          end 
        end
        control_matmul_23_8: begin
          if(_maxi_read_req_idle) begin
            control_matmul_23 <= control_matmul_23_9;
          end 
        end
        control_matmul_23_9: begin
          if(_maxi_read_idle) begin
            control_matmul_23 <= control_matmul_23_10;
          end 
        end
        control_matmul_23_10: begin
          control_matmul_23 <= control_matmul_23_11;
        end
        control_matmul_23_11: begin
          if(cparam_matmul_23_data_stationary == 0) begin
            control_matmul_23 <= control_matmul_23_12;
          end 
          if(cparam_matmul_23_data_stationary == 1) begin
            control_matmul_23 <= control_matmul_23_18;
          end 
        end
        control_matmul_23_12: begin
          control_matmul_23 <= control_matmul_23_13;
          if(matmul_23_skip_read_act) begin
            control_matmul_23 <= control_matmul_23_17;
          end 
        end
        control_matmul_23_13: begin
          control_matmul_23 <= control_matmul_23_14;
          if(matmul_23_mux_dma_pad_mask_0 || !matmul_23_mux_dma_flag_0) begin
            control_matmul_23 <= control_matmul_23_16;
          end 
        end
        control_matmul_23_14: begin
          if(_maxi_read_req_idle) begin
            control_matmul_23 <= control_matmul_23_15;
          end 
        end
        control_matmul_23_15: begin
          if(_maxi_read_idle) begin
            control_matmul_23 <= control_matmul_23_16;
          end 
        end
        control_matmul_23_16: begin
          control_matmul_23 <= control_matmul_23_17;
        end
        control_matmul_23_17: begin
          if(cparam_matmul_23_data_stationary == 0) begin
            control_matmul_23 <= control_matmul_23_18;
          end 
          if(cparam_matmul_23_data_stationary == 1) begin
            control_matmul_23 <= control_matmul_23_7;
          end 
        end
        control_matmul_23_18: begin
          if(_maxi_write_idle) begin
            control_matmul_23 <= control_matmul_23_19;
          end 
        end
        control_matmul_23_19: begin
          if(matmul_23_comp_fsm == 0) begin
            control_matmul_23 <= control_matmul_23_20;
          end 
        end
        control_matmul_23_20: begin
          control_matmul_23 <= control_matmul_23_21;
          if(matmul_23_skip_write_out) begin
            control_matmul_23 <= control_matmul_23_26;
          end 
          if((cparam_matmul_23_data_stationary == 1) && (matmul_23_prev_och_count < cparam_matmul_23_max_och_count)) begin
            control_matmul_23 <= control_matmul_23_26;
          end 
        end
        control_matmul_23_21: begin
          if(matmul_23_sync_comp_count >= matmul_23_sync_out_count + cparam_matmul_23_inc_sync_out) begin
            control_matmul_23 <= control_matmul_23_22;
          end 
        end
        control_matmul_23_22: begin
          if(!matmul_23_dma_out_mask_0) begin
            control_matmul_23 <= control_matmul_23_23;
          end 
          if(matmul_23_dma_out_mask_0) begin
            control_matmul_23 <= control_matmul_23_24;
          end 
        end
        control_matmul_23_23: begin
          if(_maxi_write_req_idle) begin
            control_matmul_23 <= control_matmul_23_24;
          end 
        end
        control_matmul_23_24: begin
          control_matmul_23 <= control_matmul_23_25;
        end
        control_matmul_23_25: begin
          matmul_23_write_count <= matmul_23_write_count + 1;
          if(matmul_23_out_ram_select == 0) begin
            matmul_23_out_laddr_offset <= matmul_23_out_laddr_offset + matmul_23_next_out_write_size;
          end 
          if((cparam_matmul_23_data_stationary == 0) && !cparam_matmul_23_keep_filter) begin
            matmul_23_out_base_offset_col <= matmul_23_out_base_offset_col + cparam_matmul_23_out_col_step;
            matmul_23_out_col_count <= matmul_23_out_col_count + 1;
          end 
          matmul_23_out_ram_select <= matmul_23_out_ram_select + 1;
          if(matmul_23_out_ram_select == 0) begin
            matmul_23_out_ram_select <= 0;
          end 
          matmul_23_sync_out_count <= matmul_23_sync_out_count + cparam_matmul_23_inc_sync_out;
          if((cparam_matmul_23_data_stationary == 0) && !cparam_matmul_23_keep_filter && (matmul_23_write_count >= cparam_matmul_23_out_num_col - 1) || (cparam_matmul_23_data_stationary == 0) && cparam_matmul_23_keep_filter || (cparam_matmul_23_data_stationary == 1)) begin
            matmul_23_sync_out_count <= matmul_23_sync_out_count + (cparam_matmul_23_inc_sync_out + cparam_matmul_23_inc_sync_out_res);
          end 
          if((cparam_matmul_23_data_stationary == 0) && !cparam_matmul_23_keep_filter) begin
            control_matmul_23 <= control_matmul_23_20;
          end 
          if((cparam_matmul_23_data_stationary == 0) && !cparam_matmul_23_keep_filter && (matmul_23_write_count >= cparam_matmul_23_out_num_col - 1) || (cparam_matmul_23_data_stationary == 0) && cparam_matmul_23_keep_filter || (cparam_matmul_23_data_stationary == 1)) begin
            control_matmul_23 <= control_matmul_23_26;
          end 
        end
        control_matmul_23_26: begin
          if(matmul_23_update_filter) begin
            matmul_23_filter_base_offset <= matmul_23_filter_base_offset + cparam_matmul_23_filter_base_step;
          end 
          if((cparam_matmul_23_data_stationary == 1) && (matmul_23_och_count >= cparam_matmul_23_max_och_count)) begin
            matmul_23_filter_base_offset <= 0;
          end 
          if(matmul_23_update_filter) begin
            matmul_23_och_count <= matmul_23_och_count + cparam_matmul_23_och_count_step;
          end 
          if((cparam_matmul_23_data_stationary == 1) && (matmul_23_och_count >= cparam_matmul_23_max_och_count)) begin
            matmul_23_och_count <= 0;
          end 
          if(matmul_23_update_filter) begin
            matmul_23_filter_page_comp_offset <= matmul_23_filter_page_comp_offset + cparam_matmul_23_filter_read_step;
            matmul_23_filter_page_dma_offset <= matmul_23_filter_page_dma_offset + cparam_matmul_23_filter_read_step;
          end 
          if(matmul_23_update_filter && (matmul_23_filter_page_comp_offset + cparam_matmul_23_filter_read_step + cparam_matmul_23_filter_read_step > 16384)) begin
            matmul_23_filter_page_comp_offset <= 0;
            matmul_23_filter_page_dma_offset <= 0;
          end 
          if(matmul_23_update_act) begin
            matmul_23_act_base_offset_row <= matmul_23_act_base_offset_row + cparam_matmul_23_act_row_step;
          end 
          if(matmul_23_update_act && (matmul_23_row_count >= cparam_matmul_23_max_row_count)) begin
            matmul_23_act_base_offset_row <= 0;
            matmul_23_act_base_offset_bat <= matmul_23_act_base_offset_bat + cparam_matmul_23_act_bat_step;
          end 
          if(matmul_23_update_act && (matmul_23_row_count >= cparam_matmul_23_max_row_count) && (matmul_23_bat_count >= cparam_matmul_23_max_bat_count)) begin
            matmul_23_act_base_offset_bat <= 0;
          end 
          if(!matmul_23_update_act) begin
            matmul_23_dma_flag_0 <= 0;
          end 
          if(matmul_23_update_act) begin
            matmul_23_dma_flag_0 <= cparam_matmul_23_dma_flag_conds_0;
          end 
          if(matmul_23_update_act && (matmul_23_row_count >= cparam_matmul_23_max_row_count)) begin
            matmul_23_dma_flag_0 <= 1;
          end 
          if(matmul_23_update_act) begin
            matmul_23_row_count <= matmul_23_row_count + cparam_matmul_23_stride_row_par_row;
          end 
          if(matmul_23_update_act && (matmul_23_row_count >= cparam_matmul_23_max_row_count)) begin
            matmul_23_row_count <= 0;
            matmul_23_bat_count <= matmul_23_bat_count + 1;
          end 
          if(matmul_23_update_act && (matmul_23_row_count >= cparam_matmul_23_max_row_count) && (matmul_23_bat_count >= cparam_matmul_23_max_bat_count)) begin
            matmul_23_bat_count <= 0;
          end 
          if(matmul_23_update_act && (cparam_matmul_23_stride_row_par_row < 1)) begin
            matmul_23_row_select <= matmul_23_row_select + cparam_matmul_23_stride_row_par_row;
            matmul_23_prev_row_select <= matmul_23_row_select;
          end 
          if(matmul_23_update_act && (cparam_matmul_23_stride_row_par_row < 1) && (matmul_23_row_select + cparam_matmul_23_stride_row_par_row >= 1)) begin
            matmul_23_row_select <= matmul_23_row_select - (1 - cparam_matmul_23_stride_row_par_row);
            matmul_23_prev_row_select <= matmul_23_row_select;
          end 
          if(matmul_23_update_act && !(cparam_matmul_23_stride_row_par_row < 1)) begin
            matmul_23_row_select <= 0;
            matmul_23_prev_row_select <= 0;
          end 
          if(matmul_23_update_act && (matmul_23_row_count >= cparam_matmul_23_max_row_count)) begin
            matmul_23_row_select <= 0;
            matmul_23_prev_row_select <= 0;
          end 
          if(matmul_23_update_act && matmul_23_mux_next_dma_flag_0) begin
            matmul_23_act_page_comp_offset_0 <= matmul_23_act_page_comp_offset_0 + cparam_matmul_23_act_read_step;
            matmul_23_act_page_dma_offset_0 <= matmul_23_act_page_dma_offset_0 + cparam_matmul_23_act_read_step;
          end 
          if(matmul_23_update_act && matmul_23_mux_next_dma_flag_0 && (matmul_23_act_page_comp_offset_0 + cparam_matmul_23_act_read_step + cparam_matmul_23_act_read_step > 4096)) begin
            matmul_23_act_page_comp_offset_0 <= 0;
            matmul_23_act_page_dma_offset_0 <= 0;
          end 
          if((cparam_matmul_23_data_stationary == 0) && (matmul_23_row_count >= cparam_matmul_23_max_row_count) && (matmul_23_bat_count >= cparam_matmul_23_max_bat_count) && cparam_matmul_23_keep_input) begin
            matmul_23_act_page_comp_offset_0 <= 0;
            matmul_23_act_page_dma_offset_0 <= 0;
          end 
          matmul_23_next_out_write_size <= (matmul_23_och_count >= cparam_matmul_23_max_och_count)? cparam_matmul_23_out_write_size_res : cparam_matmul_23_out_write_size;
          if(!matmul_23_skip_write_out) begin
            matmul_23_write_count <= 0;
            matmul_23_out_laddr_offset <= 0;
            matmul_23_out_ram_select <= 0;
          end 
          if((cparam_matmul_23_data_stationary == 0) && !matmul_23_skip_write_out) begin
            matmul_23_out_base_offset_col <= 0;
            matmul_23_out_base_offset_row <= matmul_23_out_base_offset_row + cparam_matmul_23_out_row_step;
            matmul_23_out_col_count <= 0;
            matmul_23_out_row_count <= matmul_23_out_row_count + 1;
          end 
          if((cparam_matmul_23_data_stationary == 0) && !matmul_23_skip_write_out && (matmul_23_prev_row_count >= cparam_matmul_23_max_row_count)) begin
            matmul_23_out_base_offset_row <= 0;
            matmul_23_out_base_offset_bat <= matmul_23_out_base_offset_bat + cparam_matmul_23_out_bat_step;
            matmul_23_out_row_count <= 0;
          end 
          if((cparam_matmul_23_data_stationary == 0) && !matmul_23_skip_write_out && (matmul_23_prev_row_count >= cparam_matmul_23_max_row_count) && (matmul_23_prev_bat_count >= cparam_matmul_23_max_bat_count)) begin
            matmul_23_out_base_offset_bat <= 0;
            matmul_23_out_base_offset_och <= matmul_23_out_base_offset_och + cparam_matmul_23_out_och_step;
          end 
          if((cparam_matmul_23_data_stationary == 1) && (matmul_23_prev_och_count >= cparam_matmul_23_max_och_count) && !matmul_23_skip_write_out) begin
            matmul_23_out_base_offset_row <= matmul_23_out_base_offset_row + cparam_matmul_23_out_row_step;
          end 
          if((cparam_matmul_23_data_stationary == 0) && !matmul_23_out_page) begin
            matmul_23_out_page_comp_offset <= 256;
            matmul_23_out_page_dma_offset <= 0;
            matmul_23_out_page <= 1;
          end 
          if((cparam_matmul_23_data_stationary == 0) && matmul_23_out_page) begin
            matmul_23_out_page_comp_offset <= 0;
            matmul_23_out_page_dma_offset <= 256;
            matmul_23_out_page <= 0;
          end 
          if((cparam_matmul_23_data_stationary == 1) && (matmul_23_och_count >= cparam_matmul_23_max_och_count) && !matmul_23_out_page) begin
            matmul_23_out_page_comp_offset <= 256;
            matmul_23_out_page_dma_offset <= 0;
            matmul_23_out_page <= 1;
          end 
          if((cparam_matmul_23_data_stationary == 1) && (matmul_23_och_count >= cparam_matmul_23_max_och_count) && matmul_23_out_page) begin
            matmul_23_out_page_comp_offset <= 0;
            matmul_23_out_page_dma_offset <= 256;
            matmul_23_out_page <= 0;
          end 
          matmul_23_prev_row_count <= matmul_23_row_count;
          matmul_23_prev_bat_count <= matmul_23_bat_count;
          matmul_23_prev_och_count <= matmul_23_och_count;
          if((matmul_23_row_count >= cparam_matmul_23_max_row_count) && (matmul_23_bat_count >= cparam_matmul_23_max_bat_count) && (matmul_23_och_count >= cparam_matmul_23_max_och_count)) begin
            matmul_23_skip_read_filter <= 1;
          end 
          if((cparam_matmul_23_data_stationary == 1) && cparam_matmul_23_keep_filter) begin
            matmul_23_skip_read_filter <= 1;
          end 
          if((matmul_23_row_count >= cparam_matmul_23_max_row_count) && (matmul_23_bat_count >= cparam_matmul_23_max_bat_count) && (matmul_23_och_count >= cparam_matmul_23_max_och_count)) begin
            matmul_23_skip_read_act <= 1;
          end 
          if((cparam_matmul_23_data_stationary == 0) && (matmul_23_row_count >= cparam_matmul_23_max_row_count) && (matmul_23_bat_count >= cparam_matmul_23_max_bat_count) && cparam_matmul_23_keep_input) begin
            matmul_23_skip_read_act <= 1;
          end 
          if((matmul_23_row_count >= cparam_matmul_23_max_row_count) && (matmul_23_bat_count >= cparam_matmul_23_max_bat_count) && (matmul_23_och_count >= cparam_matmul_23_max_och_count)) begin
            matmul_23_skip_comp <= 1;
          end 
          if(matmul_23_skip_write_out && (matmul_23_prev_row_count == 0) && (matmul_23_prev_bat_count == 0) && (matmul_23_prev_och_count == 0)) begin
            matmul_23_skip_write_out <= 0;
          end 
          if(cparam_matmul_23_data_stationary == 0) begin
            control_matmul_23 <= control_matmul_23_12;
          end 
          if((cparam_matmul_23_data_stationary == 0) && (matmul_23_row_count >= cparam_matmul_23_max_row_count) && (matmul_23_bat_count >= cparam_matmul_23_max_bat_count)) begin
            control_matmul_23 <= control_matmul_23_7;
          end 
          if(cparam_matmul_23_data_stationary == 1) begin
            control_matmul_23 <= control_matmul_23_7;
          end 
          if((cparam_matmul_23_data_stationary == 1) && (matmul_23_och_count >= cparam_matmul_23_max_och_count)) begin
            control_matmul_23 <= control_matmul_23_12;
          end 
          if(!matmul_23_skip_write_out && (matmul_23_prev_och_count >= cparam_matmul_23_max_och_count) && (matmul_23_prev_row_count >= cparam_matmul_23_max_row_count) && (matmul_23_prev_bat_count >= cparam_matmul_23_max_bat_count)) begin
            control_matmul_23 <= control_matmul_23_27;
          end 
        end
        control_matmul_23_27: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_matmul_23 <= control_matmul_23_28;
          end 
        end
        control_matmul_23_28: begin
          if(main_fsm == 67) begin
            _control_matmul_23_called <= 0;
          end 
          if(main_fsm == 77) begin
            _control_matmul_23_called <= 0;
          end 
          if(main_fsm == 67) begin
            control_matmul_23 <= control_matmul_23_init;
          end 
          if(main_fsm == 77) begin
            control_matmul_23 <= control_matmul_23_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_27_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_27 <= write_burst_packed_fsm_27_init;
      write_burst_packed_addr_1311 <= 0;
      write_burst_packed_stride_1312 <= 0;
      write_burst_packed_length_1313 <= 0;
      write_burst_packed_done_1314 <= 0;
    end else begin
      case(write_burst_packed_fsm_27)
        write_burst_packed_fsm_27_init: begin
          write_burst_packed_addr_1311 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_1312 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_1313 <= _maxi_read_local_size_buf;
          write_burst_packed_done_1314 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 8) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_27 <= write_burst_packed_fsm_27_1;
          end 
        end
        write_burst_packed_fsm_27_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_1311 <= write_burst_packed_addr_1311 + write_burst_packed_stride_1312;
            write_burst_packed_length_1313 <= write_burst_packed_length_1313 - 1;
            write_burst_packed_done_1314 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1313 <= 1)) begin
            write_burst_packed_done_1314 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_1314 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1313 <= 1)) begin
            write_burst_packed_fsm_27 <= write_burst_packed_fsm_27_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_27 <= write_burst_packed_fsm_27_init;
          end 
          if(0) begin
            write_burst_packed_fsm_27 <= write_burst_packed_fsm_27_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_28_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_28 <= write_burst_packed_fsm_28_init;
      write_burst_packed_addr_1324 <= 0;
      write_burst_packed_stride_1325 <= 0;
      write_burst_packed_length_1326 <= 0;
      write_burst_packed_done_1327 <= 0;
    end else begin
      case(write_burst_packed_fsm_28)
        write_burst_packed_fsm_28_init: begin
          write_burst_packed_addr_1324 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_1325 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_1326 <= _maxi_read_local_size_buf;
          write_burst_packed_done_1327 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 9) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_28 <= write_burst_packed_fsm_28_1;
          end 
        end
        write_burst_packed_fsm_28_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_1324 <= write_burst_packed_addr_1324 + write_burst_packed_stride_1325;
            write_burst_packed_length_1326 <= write_burst_packed_length_1326 - 1;
            write_burst_packed_done_1327 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1326 <= 1)) begin
            write_burst_packed_done_1327 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_1327 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1326 <= 1)) begin
            write_burst_packed_fsm_28 <= write_burst_packed_fsm_28_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_28 <= write_burst_packed_fsm_28_init;
          end 
          if(0) begin
            write_burst_packed_fsm_28 <= write_burst_packed_fsm_28_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_29_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_29 <= write_burst_packed_fsm_29_init;
      write_burst_packed_addr_1337 <= 0;
      write_burst_packed_stride_1338 <= 0;
      write_burst_packed_length_1339 <= 0;
      write_burst_packed_done_1340 <= 0;
    end else begin
      case(write_burst_packed_fsm_29)
        write_burst_packed_fsm_29_init: begin
          write_burst_packed_addr_1337 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_1338 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_1339 <= _maxi_read_local_size_buf;
          write_burst_packed_done_1340 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 10) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_29 <= write_burst_packed_fsm_29_1;
          end 
        end
        write_burst_packed_fsm_29_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_1337 <= write_burst_packed_addr_1337 + write_burst_packed_stride_1338;
            write_burst_packed_length_1339 <= write_burst_packed_length_1339 - 1;
            write_burst_packed_done_1340 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1339 <= 1)) begin
            write_burst_packed_done_1340 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_1340 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1339 <= 1)) begin
            write_burst_packed_fsm_29 <= write_burst_packed_fsm_29_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_29 <= write_burst_packed_fsm_29_init;
          end 
          if(0) begin
            write_burst_packed_fsm_29 <= write_burst_packed_fsm_29_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_30_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_30 <= write_burst_packed_fsm_30_init;
      write_burst_packed_addr_1350 <= 0;
      write_burst_packed_stride_1351 <= 0;
      write_burst_packed_length_1352 <= 0;
      write_burst_packed_done_1353 <= 0;
    end else begin
      case(write_burst_packed_fsm_30)
        write_burst_packed_fsm_30_init: begin
          write_burst_packed_addr_1350 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_1351 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_1352 <= _maxi_read_local_size_buf;
          write_burst_packed_done_1353 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 11) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_30 <= write_burst_packed_fsm_30_1;
          end 
        end
        write_burst_packed_fsm_30_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_1350 <= write_burst_packed_addr_1350 + write_burst_packed_stride_1351;
            write_burst_packed_length_1352 <= write_burst_packed_length_1352 - 1;
            write_burst_packed_done_1353 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1352 <= 1)) begin
            write_burst_packed_done_1353 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_1353 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1352 <= 1)) begin
            write_burst_packed_fsm_30 <= write_burst_packed_fsm_30_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_30 <= write_burst_packed_fsm_30_init;
          end 
          if(0) begin
            write_burst_packed_fsm_30 <= write_burst_packed_fsm_30_init;
          end 
        end
      endcase
    end
  end

  localparam matmul_23_comp_fsm_1 = 1;
  localparam matmul_23_comp_fsm_2 = 2;
  localparam matmul_23_comp_fsm_3 = 3;
  localparam matmul_23_comp_fsm_4 = 4;
  localparam matmul_23_comp_fsm_5 = 5;
  localparam matmul_23_comp_fsm_6 = 6;

  always @(posedge CLK) begin
    if(RST) begin
      matmul_23_comp_fsm <= matmul_23_comp_fsm_init;
      matmul_23_stream_act_local_0 <= 0;
      matmul_23_stream_out_local_col <= 0;
      matmul_23_stream_out_local_val <= 0;
      matmul_23_col_count <= 0;
      matmul_23_col_select <= 0;
      matmul_23_filter_page_comp_offset_buf <= 0;
      matmul_23_act_page_comp_offset_buf_0 <= 0;
      matmul_23_out_page_comp_offset_buf <= 0;
      matmul_23_row_count_buf <= 0;
      matmul_23_row_select_buf <= 0;
      matmul_23_och_count_buf <= 0;
      matmul_23_next_stream_num_ops <= 0;
      matmul_23_stream_pad_masks <= 0;
      matmul_23_sync_comp_count <= 0;
    end else begin
      if(_stream_matmul_23_sink_stop) begin
        matmul_23_sync_comp_count <= matmul_23_sync_comp_count + 1;
      end 
      if(control_matmul_23 == 6) begin
        matmul_23_sync_comp_count <= 0;
      end 
      case(matmul_23_comp_fsm)
        matmul_23_comp_fsm_init: begin
          if((control_matmul_23 == 19) && !matmul_23_skip_comp) begin
            matmul_23_comp_fsm <= matmul_23_comp_fsm_1;
          end 
        end
        matmul_23_comp_fsm_1: begin
          matmul_23_stream_act_local_0 <= 0;
          if(cparam_matmul_23_stream_act_local_small_flags_0) begin
            matmul_23_stream_act_local_0 <= cparam_matmul_23_stream_act_local_small_offset;
          end 
          if(cparam_matmul_23_stream_act_local_large_flags_0) begin
            matmul_23_stream_act_local_0 <= cparam_matmul_23_stream_act_local_large_offset;
          end 
          matmul_23_stream_out_local_col <= 0;
          if((cparam_matmul_23_data_stationary == 1) && (matmul_23_och_count == 0)) begin
            matmul_23_stream_out_local_val <= 0;
          end 
          matmul_23_col_count <= 0;
          matmul_23_col_select <= cparam_matmul_23_col_select_initval;
          matmul_23_filter_page_comp_offset_buf <= matmul_23_filter_page_comp_offset;
          matmul_23_act_page_comp_offset_buf_0 <= matmul_23_act_page_comp_offset_0;
          matmul_23_out_page_comp_offset_buf <= matmul_23_out_page_comp_offset;
          matmul_23_row_count_buf <= matmul_23_row_count;
          matmul_23_row_select_buf <= matmul_23_row_select;
          matmul_23_och_count_buf <= matmul_23_och_count;
          matmul_23_next_stream_num_ops <= (matmul_23_och_count >= cparam_matmul_23_max_och_count)? cparam_matmul_23_stream_num_ops_res : cparam_matmul_23_stream_num_ops;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_2;
        end
        matmul_23_comp_fsm_2: begin
          matmul_23_stream_pad_masks <= { matmul_23_stream_pad_mask_0_0 };
          matmul_23_comp_fsm <= matmul_23_comp_fsm_3;
        end
        matmul_23_comp_fsm_3: begin
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          if(_stream_matmul_23_stream_oready) begin
            matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
          end 
          matmul_23_comp_fsm <= matmul_23_comp_fsm_4;
        end
        matmul_23_comp_fsm_4: begin
          if(!_stream_matmul_23_source_busy) begin
            matmul_23_comp_fsm <= matmul_23_comp_fsm_5;
          end 
        end
        matmul_23_comp_fsm_5: begin
          if(_stream_matmul_23_busy) begin
            matmul_23_comp_fsm <= matmul_23_comp_fsm_6;
          end 
        end
        matmul_23_comp_fsm_6: begin
          if(!((matmul_23_col_select == 0)? cparam_matmul_23_inc_act_laddr_conds_0 : 0)) begin
            matmul_23_stream_act_local_0 <= matmul_23_stream_act_local_0 + cparam_matmul_23_inc_act_laddr_small;
          end 
          if((matmul_23_col_select == 0)? cparam_matmul_23_inc_act_laddr_conds_0 : 0) begin
            matmul_23_stream_act_local_0 <= matmul_23_stream_act_local_0 + cparam_matmul_23_inc_act_laddr_large;
          end 
          if(matmul_23_col_count >= cparam_matmul_23_max_col_count) begin
            matmul_23_stream_act_local_0 <= 0;
          end 
          if((matmul_23_col_count >= cparam_matmul_23_max_col_count) && cparam_matmul_23_stream_act_local_small_flags_0) begin
            matmul_23_stream_act_local_0 <= cparam_matmul_23_stream_act_local_small_offset;
          end 
          if((matmul_23_col_count >= cparam_matmul_23_max_col_count) && cparam_matmul_23_stream_act_local_large_flags_0) begin
            matmul_23_stream_act_local_0 <= cparam_matmul_23_stream_act_local_large_offset;
          end 
          if(cparam_matmul_23_data_stationary == 0) begin
            matmul_23_stream_out_local_col <= matmul_23_stream_out_local_col + matmul_23_next_stream_num_ops;
          end 
          if((cparam_matmul_23_data_stationary == 0) && (matmul_23_col_count >= cparam_matmul_23_max_col_count)) begin
            matmul_23_stream_out_local_col <= 0;
          end 
          if(cparam_matmul_23_data_stationary == 1) begin
            matmul_23_stream_out_local_col <= matmul_23_stream_out_local_col + cparam_matmul_23_inc_out_laddr_col;
          end 
          if((cparam_matmul_23_data_stationary == 1) && (matmul_23_col_count >= cparam_matmul_23_max_col_count)) begin
            matmul_23_stream_out_local_val <= matmul_23_stream_out_local_val + matmul_23_next_stream_num_ops;
            matmul_23_stream_out_local_col <= 0;
          end 
          matmul_23_col_count <= matmul_23_col_count + cparam_matmul_23_stride_col_par_col;
          if(matmul_23_col_count >= cparam_matmul_23_max_col_count) begin
            matmul_23_col_count <= 0;
          end 
          matmul_23_col_select <= matmul_23_col_select + cparam_matmul_23_stride_col_mod_filter_num;
          if(matmul_23_col_select + cparam_matmul_23_stride_col_mod_filter_num >= 1) begin
            matmul_23_col_select <= matmul_23_col_select - cparam_matmul_23_filter_num_col_minus_stride_col_mod;
          end 
          if(matmul_23_col_count >= cparam_matmul_23_max_col_count) begin
            matmul_23_col_select <= cparam_matmul_23_col_select_initval;
          end 
          matmul_23_comp_fsm <= matmul_23_comp_fsm_2;
          if(matmul_23_col_count >= cparam_matmul_23_max_col_count) begin
            matmul_23_comp_fsm <= matmul_23_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_23_source_7_source_pat_fsm_0_1 = 1;
  localparam _stream_matmul_23_source_7_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_23_source_7_source_pat_fsm_0 <= _stream_matmul_23_source_7_source_pat_fsm_0_init;
    end else begin
      case(_stream_matmul_23_source_7_source_pat_fsm_0)
        _stream_matmul_23_source_7_source_pat_fsm_0_init: begin
          if(_stream_matmul_23_source_start && _stream_matmul_23_source_7_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_7_source_pat_fsm_0 <= _stream_matmul_23_source_7_source_pat_fsm_0_1;
          end 
        end
        _stream_matmul_23_source_7_source_pat_fsm_0_1: begin
          if(_stream_matmul_23_source_stop && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_7_source_pat_fsm_0 <= _stream_matmul_23_source_7_source_pat_fsm_0_init;
          end 
          if((_source_stream_matmul_23_source_7_pat_count_0 == 0) && (_source_stream_matmul_23_source_7_pat_count_1 == 0) && (_source_stream_matmul_23_source_7_pat_count_2 == 0) && (_source_stream_matmul_23_source_7_pat_count_3 == 0) && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_7_source_pat_fsm_0 <= _stream_matmul_23_source_7_source_pat_fsm_0_2;
          end 
        end
        _stream_matmul_23_source_7_source_pat_fsm_0_2: begin
          if(_stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_7_source_pat_fsm_0 <= _stream_matmul_23_source_7_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_23_source_9_source_pat_fsm_1_1 = 1;
  localparam _stream_matmul_23_source_9_source_pat_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_23_source_9_source_pat_fsm_1 <= _stream_matmul_23_source_9_source_pat_fsm_1_init;
    end else begin
      case(_stream_matmul_23_source_9_source_pat_fsm_1)
        _stream_matmul_23_source_9_source_pat_fsm_1_init: begin
          if(_stream_matmul_23_source_start && _stream_matmul_23_source_9_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_9_source_pat_fsm_1 <= _stream_matmul_23_source_9_source_pat_fsm_1_1;
          end 
        end
        _stream_matmul_23_source_9_source_pat_fsm_1_1: begin
          if(_stream_matmul_23_source_stop && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_9_source_pat_fsm_1 <= _stream_matmul_23_source_9_source_pat_fsm_1_init;
          end 
          if((_source_stream_matmul_23_source_9_pat_count_0 == 0) && (_source_stream_matmul_23_source_9_pat_count_1 == 0) && (_source_stream_matmul_23_source_9_pat_count_2 == 0) && (_source_stream_matmul_23_source_9_pat_count_3 == 0) && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_9_source_pat_fsm_1 <= _stream_matmul_23_source_9_source_pat_fsm_1_2;
          end 
        end
        _stream_matmul_23_source_9_source_pat_fsm_1_2: begin
          if(_stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_9_source_pat_fsm_1 <= _stream_matmul_23_source_9_source_pat_fsm_1_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_1395 <= 0;
    end else begin
      if(_stream_matmul_23_stream_oready && _stream_matmul_23_source_20_source_ram_renable && (_stream_matmul_23_source_20_source_sel == 3)) begin
        _tmp_1395 <= read_rtl_bank_1394;
      end 
    end
  end

  localparam _stream_matmul_23_source_20_source_pat_fsm_2_1 = 1;
  localparam _stream_matmul_23_source_20_source_pat_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_23_source_20_source_pat_fsm_2 <= _stream_matmul_23_source_20_source_pat_fsm_2_init;
    end else begin
      case(_stream_matmul_23_source_20_source_pat_fsm_2)
        _stream_matmul_23_source_20_source_pat_fsm_2_init: begin
          if(_stream_matmul_23_source_start && _stream_matmul_23_source_20_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_20_source_pat_fsm_2 <= _stream_matmul_23_source_20_source_pat_fsm_2_1;
          end 
        end
        _stream_matmul_23_source_20_source_pat_fsm_2_1: begin
          if(_stream_matmul_23_source_stop && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_20_source_pat_fsm_2 <= _stream_matmul_23_source_20_source_pat_fsm_2_init;
          end 
          if((_source_stream_matmul_23_source_20_pat_count_0 == 0) && (_source_stream_matmul_23_source_20_pat_count_1 == 0) && (_source_stream_matmul_23_source_20_pat_count_2 == 0) && (_source_stream_matmul_23_source_20_pat_count_3 == 0) && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_20_source_pat_fsm_2 <= _stream_matmul_23_source_20_source_pat_fsm_2_2;
          end 
        end
        _stream_matmul_23_source_20_source_pat_fsm_2_2: begin
          if(_stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_20_source_pat_fsm_2 <= _stream_matmul_23_source_20_source_pat_fsm_2_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_1404 <= 0;
    end else begin
      if(_stream_matmul_23_stream_oready && _stream_matmul_23_source_21_source_ram_renable && (_stream_matmul_23_source_21_source_sel == 4)) begin
        _tmp_1404 <= read_rtl_bank_1403;
      end 
    end
  end

  localparam _stream_matmul_23_source_21_source_pat_fsm_3_1 = 1;
  localparam _stream_matmul_23_source_21_source_pat_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_23_source_21_source_pat_fsm_3 <= _stream_matmul_23_source_21_source_pat_fsm_3_init;
    end else begin
      case(_stream_matmul_23_source_21_source_pat_fsm_3)
        _stream_matmul_23_source_21_source_pat_fsm_3_init: begin
          if(_stream_matmul_23_source_start && _stream_matmul_23_source_21_source_mode & 5'b10 && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_21_source_pat_fsm_3 <= _stream_matmul_23_source_21_source_pat_fsm_3_1;
          end 
        end
        _stream_matmul_23_source_21_source_pat_fsm_3_1: begin
          if(_stream_matmul_23_source_stop && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_21_source_pat_fsm_3 <= _stream_matmul_23_source_21_source_pat_fsm_3_init;
          end 
          if((_source_stream_matmul_23_source_21_pat_count_0 == 0) && (_source_stream_matmul_23_source_21_pat_count_1 == 0) && (_source_stream_matmul_23_source_21_pat_count_2 == 0) && (_source_stream_matmul_23_source_21_pat_count_3 == 0) && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_21_source_pat_fsm_3 <= _stream_matmul_23_source_21_source_pat_fsm_3_2;
          end 
        end
        _stream_matmul_23_source_21_source_pat_fsm_3_2: begin
          if(_stream_matmul_23_stream_oready) begin
            _stream_matmul_23_source_21_source_pat_fsm_3 <= _stream_matmul_23_source_21_source_pat_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_23_sink_26_sink_fsm_4_1 = 1;
  localparam _stream_matmul_23_sink_26_sink_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_23_sink_26_sink_fsm_4 <= _stream_matmul_23_sink_26_sink_fsm_4_init;
    end else begin
      case(_stream_matmul_23_sink_26_sink_fsm_4)
        _stream_matmul_23_sink_26_sink_fsm_4_init: begin
          if(_stream_matmul_23_sink_start && _stream_matmul_23_sink_26_sink_mode & 5'b1 && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_sink_26_sink_fsm_4 <= _stream_matmul_23_sink_26_sink_fsm_4_1;
          end 
        end
        _stream_matmul_23_sink_26_sink_fsm_4_1: begin
          if(_stream_matmul_23_stream_oready) begin
            _stream_matmul_23_sink_26_sink_fsm_4 <= _stream_matmul_23_sink_26_sink_fsm_4_2;
          end 
        end
        _stream_matmul_23_sink_26_sink_fsm_4_2: begin
          if(stream_matmul_23_sink_27_data && (_stream_matmul_23_sink_26_sink_count == 1) && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_sink_26_sink_fsm_4 <= _stream_matmul_23_sink_26_sink_fsm_4_init;
          end 
          if(_stream_matmul_23_sink_stop && _stream_matmul_23_stream_oready) begin
            _stream_matmul_23_sink_26_sink_fsm_4 <= _stream_matmul_23_sink_26_sink_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam control_matmul_33_1 = 1;
  localparam control_matmul_33_2 = 2;
  localparam control_matmul_33_3 = 3;
  localparam control_matmul_33_4 = 4;
  localparam control_matmul_33_5 = 5;
  localparam control_matmul_33_6 = 6;
  localparam control_matmul_33_7 = 7;
  localparam control_matmul_33_8 = 8;
  localparam control_matmul_33_9 = 9;
  localparam control_matmul_33_10 = 10;
  localparam control_matmul_33_11 = 11;
  localparam control_matmul_33_12 = 12;
  localparam control_matmul_33_13 = 13;
  localparam control_matmul_33_14 = 14;
  localparam control_matmul_33_15 = 15;
  localparam control_matmul_33_16 = 16;
  localparam control_matmul_33_17 = 17;
  localparam control_matmul_33_18 = 18;
  localparam control_matmul_33_19 = 19;
  localparam control_matmul_33_20 = 20;
  localparam control_matmul_33_21 = 21;
  localparam control_matmul_33_22 = 22;
  localparam control_matmul_33_23 = 23;
  localparam control_matmul_33_24 = 24;
  localparam control_matmul_33_25 = 25;
  localparam control_matmul_33_26 = 26;
  localparam control_matmul_33_27 = 27;
  localparam control_matmul_33_28 = 28;

  always @(posedge CLK) begin
    if(RST) begin
      control_matmul_33 <= control_matmul_33_init;
      _control_matmul_33_called <= 0;
      matmul_33_filter_base_offset <= 0;
      matmul_33_filter_page_comp_offset <= 0;
      matmul_33_filter_page_dma_offset <= 0;
      matmul_33_act_base_offset_row <= 0;
      matmul_33_act_base_offset_bat <= 0;
      matmul_33_dma_flag_0 <= 0;
      matmul_33_act_page_comp_offset_0 <= 0;
      matmul_33_act_page_dma_offset_0 <= 0;
      matmul_33_out_base_offset_val <= 0;
      matmul_33_out_base_offset_col <= 0;
      matmul_33_out_base_offset_row <= 0;
      matmul_33_out_base_offset_bat <= 0;
      matmul_33_out_base_offset_och <= 0;
      matmul_33_out_page <= 0;
      matmul_33_out_page_comp_offset <= 0;
      matmul_33_out_page_dma_offset <= 0;
      matmul_33_out_laddr_offset <= 0;
      matmul_33_sync_out_count <= 0;
      matmul_33_write_count <= 0;
      matmul_33_next_out_write_size <= 0;
      matmul_33_row_count <= 0;
      matmul_33_bat_count <= 0;
      matmul_33_och_count <= 0;
      matmul_33_row_select <= 0;
      matmul_33_prev_row_count <= 0;
      matmul_33_prev_bat_count <= 0;
      matmul_33_prev_och_count <= 0;
      matmul_33_prev_row_select <= 0;
      matmul_33_out_col_count <= 0;
      matmul_33_out_row_count <= 0;
      matmul_33_out_ram_select <= 0;
      matmul_33_skip_read_filter <= 0;
      matmul_33_skip_read_act <= 0;
      matmul_33_skip_comp <= 0;
      matmul_33_skip_write_out <= 1;
    end else begin
      case(control_matmul_33)
        control_matmul_33_init: begin
          if(main_fsm == 83) begin
            _control_matmul_33_called <= 1;
          end 
          if(main_fsm == 83) begin
            control_matmul_33 <= control_matmul_33_1;
          end 
        end
        control_matmul_33_1: begin
          control_matmul_33 <= control_matmul_33_2;
        end
        control_matmul_33_2: begin
          matmul_33_filter_base_offset <= 0;
          matmul_33_filter_page_comp_offset <= 0;
          matmul_33_filter_page_dma_offset <= 0;
          matmul_33_act_base_offset_row <= 0;
          matmul_33_act_base_offset_bat <= 0;
          matmul_33_dma_flag_0 <= 1;
          matmul_33_act_page_comp_offset_0 <= 0;
          matmul_33_act_page_dma_offset_0 <= 0;
          matmul_33_out_base_offset_val <= 0;
          matmul_33_out_base_offset_col <= 0;
          matmul_33_out_base_offset_row <= 0;
          matmul_33_out_base_offset_bat <= 0;
          matmul_33_out_base_offset_och <= 0;
          matmul_33_out_page <= 0;
          matmul_33_out_page_comp_offset <= 0;
          matmul_33_out_page_dma_offset <= 0;
          matmul_33_out_laddr_offset <= 0;
          matmul_33_sync_out_count <= 0;
          matmul_33_write_count <= 0;
          matmul_33_next_out_write_size <= (cparam_matmul_33_max_och_count == 0)? cparam_matmul_33_out_write_size_res : cparam_matmul_33_out_write_size;
          matmul_33_row_count <= 0;
          matmul_33_bat_count <= 0;
          matmul_33_och_count <= 0;
          matmul_33_row_select <= 0;
          matmul_33_prev_row_count <= 0;
          matmul_33_prev_bat_count <= 0;
          matmul_33_prev_och_count <= 0;
          matmul_33_prev_row_select <= 0;
          matmul_33_out_col_count <= 0;
          matmul_33_out_row_count <= 0;
          matmul_33_out_ram_select <= 0;
          matmul_33_skip_read_filter <= 0;
          matmul_33_skip_read_act <= 0;
          matmul_33_skip_comp <= 0;
          matmul_33_skip_write_out <= 1;
          if(_maxi_read_req_idle) begin
            control_matmul_33 <= control_matmul_33_3;
          end 
        end
        control_matmul_33_3: begin
          if(_maxi_read_idle) begin
            control_matmul_33 <= control_matmul_33_4;
          end 
        end
        control_matmul_33_4: begin
          if(_maxi_read_req_idle) begin
            control_matmul_33 <= control_matmul_33_5;
          end 
        end
        control_matmul_33_5: begin
          if(_maxi_read_idle) begin
            control_matmul_33 <= control_matmul_33_6;
          end 
        end
        control_matmul_33_6: begin
          if(cparam_matmul_33_data_stationary == 0) begin
            control_matmul_33 <= control_matmul_33_7;
          end 
          if(cparam_matmul_33_data_stationary == 1) begin
            control_matmul_33 <= control_matmul_33_12;
          end 
        end
        control_matmul_33_7: begin
          control_matmul_33 <= control_matmul_33_8;
          if(matmul_33_skip_read_filter) begin
            control_matmul_33 <= control_matmul_33_11;
          end 
        end
        control_matmul_33_8: begin
          if(_maxi_read_req_idle) begin
            control_matmul_33 <= control_matmul_33_9;
          end 
        end
        control_matmul_33_9: begin
          if(_maxi_read_idle) begin
            control_matmul_33 <= control_matmul_33_10;
          end 
        end
        control_matmul_33_10: begin
          control_matmul_33 <= control_matmul_33_11;
        end
        control_matmul_33_11: begin
          if(cparam_matmul_33_data_stationary == 0) begin
            control_matmul_33 <= control_matmul_33_12;
          end 
          if(cparam_matmul_33_data_stationary == 1) begin
            control_matmul_33 <= control_matmul_33_18;
          end 
        end
        control_matmul_33_12: begin
          control_matmul_33 <= control_matmul_33_13;
          if(matmul_33_skip_read_act) begin
            control_matmul_33 <= control_matmul_33_17;
          end 
        end
        control_matmul_33_13: begin
          control_matmul_33 <= control_matmul_33_14;
          if(matmul_33_mux_dma_pad_mask_0 || !matmul_33_mux_dma_flag_0) begin
            control_matmul_33 <= control_matmul_33_16;
          end 
        end
        control_matmul_33_14: begin
          if(_maxi_read_req_idle) begin
            control_matmul_33 <= control_matmul_33_15;
          end 
        end
        control_matmul_33_15: begin
          if(_maxi_read_idle) begin
            control_matmul_33 <= control_matmul_33_16;
          end 
        end
        control_matmul_33_16: begin
          control_matmul_33 <= control_matmul_33_17;
        end
        control_matmul_33_17: begin
          if(cparam_matmul_33_data_stationary == 0) begin
            control_matmul_33 <= control_matmul_33_18;
          end 
          if(cparam_matmul_33_data_stationary == 1) begin
            control_matmul_33 <= control_matmul_33_7;
          end 
        end
        control_matmul_33_18: begin
          if(_maxi_write_idle) begin
            control_matmul_33 <= control_matmul_33_19;
          end 
        end
        control_matmul_33_19: begin
          if(matmul_33_comp_fsm == 0) begin
            control_matmul_33 <= control_matmul_33_20;
          end 
        end
        control_matmul_33_20: begin
          control_matmul_33 <= control_matmul_33_21;
          if(matmul_33_skip_write_out) begin
            control_matmul_33 <= control_matmul_33_26;
          end 
          if((cparam_matmul_33_data_stationary == 1) && (matmul_33_prev_och_count < cparam_matmul_33_max_och_count)) begin
            control_matmul_33 <= control_matmul_33_26;
          end 
        end
        control_matmul_33_21: begin
          if(matmul_33_sync_comp_count >= matmul_33_sync_out_count + cparam_matmul_33_inc_sync_out) begin
            control_matmul_33 <= control_matmul_33_22;
          end 
        end
        control_matmul_33_22: begin
          if(!matmul_33_dma_out_mask_0) begin
            control_matmul_33 <= control_matmul_33_23;
          end 
          if(matmul_33_dma_out_mask_0) begin
            control_matmul_33 <= control_matmul_33_24;
          end 
        end
        control_matmul_33_23: begin
          if(_maxi_write_req_idle) begin
            control_matmul_33 <= control_matmul_33_24;
          end 
        end
        control_matmul_33_24: begin
          control_matmul_33 <= control_matmul_33_25;
        end
        control_matmul_33_25: begin
          matmul_33_write_count <= matmul_33_write_count + 1;
          if(matmul_33_out_ram_select == 0) begin
            matmul_33_out_laddr_offset <= matmul_33_out_laddr_offset + matmul_33_next_out_write_size;
          end 
          if((cparam_matmul_33_data_stationary == 0) && !cparam_matmul_33_keep_filter) begin
            matmul_33_out_base_offset_col <= matmul_33_out_base_offset_col + cparam_matmul_33_out_col_step;
            matmul_33_out_col_count <= matmul_33_out_col_count + 1;
          end 
          matmul_33_out_ram_select <= matmul_33_out_ram_select + 1;
          if(matmul_33_out_ram_select == 0) begin
            matmul_33_out_ram_select <= 0;
          end 
          matmul_33_sync_out_count <= matmul_33_sync_out_count + cparam_matmul_33_inc_sync_out;
          if((cparam_matmul_33_data_stationary == 0) && !cparam_matmul_33_keep_filter && (matmul_33_write_count >= cparam_matmul_33_out_num_col - 1) || (cparam_matmul_33_data_stationary == 0) && cparam_matmul_33_keep_filter || (cparam_matmul_33_data_stationary == 1)) begin
            matmul_33_sync_out_count <= matmul_33_sync_out_count + (cparam_matmul_33_inc_sync_out + cparam_matmul_33_inc_sync_out_res);
          end 
          if((cparam_matmul_33_data_stationary == 0) && !cparam_matmul_33_keep_filter) begin
            control_matmul_33 <= control_matmul_33_20;
          end 
          if((cparam_matmul_33_data_stationary == 0) && !cparam_matmul_33_keep_filter && (matmul_33_write_count >= cparam_matmul_33_out_num_col - 1) || (cparam_matmul_33_data_stationary == 0) && cparam_matmul_33_keep_filter || (cparam_matmul_33_data_stationary == 1)) begin
            control_matmul_33 <= control_matmul_33_26;
          end 
        end
        control_matmul_33_26: begin
          if(matmul_33_update_filter) begin
            matmul_33_filter_base_offset <= matmul_33_filter_base_offset + cparam_matmul_33_filter_base_step;
          end 
          if((cparam_matmul_33_data_stationary == 1) && (matmul_33_och_count >= cparam_matmul_33_max_och_count)) begin
            matmul_33_filter_base_offset <= 0;
          end 
          if(matmul_33_update_filter) begin
            matmul_33_och_count <= matmul_33_och_count + cparam_matmul_33_och_count_step;
          end 
          if((cparam_matmul_33_data_stationary == 1) && (matmul_33_och_count >= cparam_matmul_33_max_och_count)) begin
            matmul_33_och_count <= 0;
          end 
          if(matmul_33_update_filter) begin
            matmul_33_filter_page_comp_offset <= matmul_33_filter_page_comp_offset + cparam_matmul_33_filter_read_step;
            matmul_33_filter_page_dma_offset <= matmul_33_filter_page_dma_offset + cparam_matmul_33_filter_read_step;
          end 
          if(matmul_33_update_filter && (matmul_33_filter_page_comp_offset + cparam_matmul_33_filter_read_step + cparam_matmul_33_filter_read_step > 512)) begin
            matmul_33_filter_page_comp_offset <= 0;
            matmul_33_filter_page_dma_offset <= 0;
          end 
          if(matmul_33_update_act) begin
            matmul_33_act_base_offset_row <= matmul_33_act_base_offset_row + cparam_matmul_33_act_row_step;
          end 
          if(matmul_33_update_act && (matmul_33_row_count >= cparam_matmul_33_max_row_count)) begin
            matmul_33_act_base_offset_row <= 0;
            matmul_33_act_base_offset_bat <= matmul_33_act_base_offset_bat + cparam_matmul_33_act_bat_step;
          end 
          if(matmul_33_update_act && (matmul_33_row_count >= cparam_matmul_33_max_row_count) && (matmul_33_bat_count >= cparam_matmul_33_max_bat_count)) begin
            matmul_33_act_base_offset_bat <= 0;
          end 
          if(!matmul_33_update_act) begin
            matmul_33_dma_flag_0 <= 0;
          end 
          if(matmul_33_update_act) begin
            matmul_33_dma_flag_0 <= cparam_matmul_33_dma_flag_conds_0;
          end 
          if(matmul_33_update_act && (matmul_33_row_count >= cparam_matmul_33_max_row_count)) begin
            matmul_33_dma_flag_0 <= 1;
          end 
          if(matmul_33_update_act) begin
            matmul_33_row_count <= matmul_33_row_count + cparam_matmul_33_stride_row_par_row;
          end 
          if(matmul_33_update_act && (matmul_33_row_count >= cparam_matmul_33_max_row_count)) begin
            matmul_33_row_count <= 0;
            matmul_33_bat_count <= matmul_33_bat_count + 1;
          end 
          if(matmul_33_update_act && (matmul_33_row_count >= cparam_matmul_33_max_row_count) && (matmul_33_bat_count >= cparam_matmul_33_max_bat_count)) begin
            matmul_33_bat_count <= 0;
          end 
          if(matmul_33_update_act && (cparam_matmul_33_stride_row_par_row < 1)) begin
            matmul_33_row_select <= matmul_33_row_select + cparam_matmul_33_stride_row_par_row;
            matmul_33_prev_row_select <= matmul_33_row_select;
          end 
          if(matmul_33_update_act && (cparam_matmul_33_stride_row_par_row < 1) && (matmul_33_row_select + cparam_matmul_33_stride_row_par_row >= 1)) begin
            matmul_33_row_select <= matmul_33_row_select - (1 - cparam_matmul_33_stride_row_par_row);
            matmul_33_prev_row_select <= matmul_33_row_select;
          end 
          if(matmul_33_update_act && !(cparam_matmul_33_stride_row_par_row < 1)) begin
            matmul_33_row_select <= 0;
            matmul_33_prev_row_select <= 0;
          end 
          if(matmul_33_update_act && (matmul_33_row_count >= cparam_matmul_33_max_row_count)) begin
            matmul_33_row_select <= 0;
            matmul_33_prev_row_select <= 0;
          end 
          if(matmul_33_update_act && matmul_33_mux_next_dma_flag_0) begin
            matmul_33_act_page_comp_offset_0 <= matmul_33_act_page_comp_offset_0 + cparam_matmul_33_act_read_step;
            matmul_33_act_page_dma_offset_0 <= matmul_33_act_page_dma_offset_0 + cparam_matmul_33_act_read_step;
          end 
          if(matmul_33_update_act && matmul_33_mux_next_dma_flag_0 && (matmul_33_act_page_comp_offset_0 + cparam_matmul_33_act_read_step + cparam_matmul_33_act_read_step > 512)) begin
            matmul_33_act_page_comp_offset_0 <= 0;
            matmul_33_act_page_dma_offset_0 <= 0;
          end 
          if((cparam_matmul_33_data_stationary == 0) && (matmul_33_row_count >= cparam_matmul_33_max_row_count) && (matmul_33_bat_count >= cparam_matmul_33_max_bat_count) && cparam_matmul_33_keep_input) begin
            matmul_33_act_page_comp_offset_0 <= 0;
            matmul_33_act_page_dma_offset_0 <= 0;
          end 
          matmul_33_next_out_write_size <= (matmul_33_och_count >= cparam_matmul_33_max_och_count)? cparam_matmul_33_out_write_size_res : cparam_matmul_33_out_write_size;
          if(!matmul_33_skip_write_out) begin
            matmul_33_write_count <= 0;
            matmul_33_out_laddr_offset <= 0;
            matmul_33_out_ram_select <= 0;
          end 
          if((cparam_matmul_33_data_stationary == 0) && !matmul_33_skip_write_out) begin
            matmul_33_out_base_offset_col <= 0;
            matmul_33_out_base_offset_row <= matmul_33_out_base_offset_row + cparam_matmul_33_out_row_step;
            matmul_33_out_col_count <= 0;
            matmul_33_out_row_count <= matmul_33_out_row_count + 1;
          end 
          if((cparam_matmul_33_data_stationary == 0) && !matmul_33_skip_write_out && (matmul_33_prev_row_count >= cparam_matmul_33_max_row_count)) begin
            matmul_33_out_base_offset_row <= 0;
            matmul_33_out_base_offset_bat <= matmul_33_out_base_offset_bat + cparam_matmul_33_out_bat_step;
            matmul_33_out_row_count <= 0;
          end 
          if((cparam_matmul_33_data_stationary == 0) && !matmul_33_skip_write_out && (matmul_33_prev_row_count >= cparam_matmul_33_max_row_count) && (matmul_33_prev_bat_count >= cparam_matmul_33_max_bat_count)) begin
            matmul_33_out_base_offset_bat <= 0;
            matmul_33_out_base_offset_och <= matmul_33_out_base_offset_och + cparam_matmul_33_out_och_step;
          end 
          if((cparam_matmul_33_data_stationary == 1) && (matmul_33_prev_och_count >= cparam_matmul_33_max_och_count) && !matmul_33_skip_write_out) begin
            matmul_33_out_base_offset_row <= matmul_33_out_base_offset_row + cparam_matmul_33_out_row_step;
          end 
          if((cparam_matmul_33_data_stationary == 0) && !matmul_33_out_page) begin
            matmul_33_out_page_comp_offset <= 64;
            matmul_33_out_page_dma_offset <= 0;
            matmul_33_out_page <= 1;
          end 
          if((cparam_matmul_33_data_stationary == 0) && matmul_33_out_page) begin
            matmul_33_out_page_comp_offset <= 0;
            matmul_33_out_page_dma_offset <= 64;
            matmul_33_out_page <= 0;
          end 
          if((cparam_matmul_33_data_stationary == 1) && (matmul_33_och_count >= cparam_matmul_33_max_och_count) && !matmul_33_out_page) begin
            matmul_33_out_page_comp_offset <= 64;
            matmul_33_out_page_dma_offset <= 0;
            matmul_33_out_page <= 1;
          end 
          if((cparam_matmul_33_data_stationary == 1) && (matmul_33_och_count >= cparam_matmul_33_max_och_count) && matmul_33_out_page) begin
            matmul_33_out_page_comp_offset <= 0;
            matmul_33_out_page_dma_offset <= 64;
            matmul_33_out_page <= 0;
          end 
          matmul_33_prev_row_count <= matmul_33_row_count;
          matmul_33_prev_bat_count <= matmul_33_bat_count;
          matmul_33_prev_och_count <= matmul_33_och_count;
          if((matmul_33_row_count >= cparam_matmul_33_max_row_count) && (matmul_33_bat_count >= cparam_matmul_33_max_bat_count) && (matmul_33_och_count >= cparam_matmul_33_max_och_count)) begin
            matmul_33_skip_read_filter <= 1;
          end 
          if((cparam_matmul_33_data_stationary == 1) && cparam_matmul_33_keep_filter) begin
            matmul_33_skip_read_filter <= 1;
          end 
          if((matmul_33_row_count >= cparam_matmul_33_max_row_count) && (matmul_33_bat_count >= cparam_matmul_33_max_bat_count) && (matmul_33_och_count >= cparam_matmul_33_max_och_count)) begin
            matmul_33_skip_read_act <= 1;
          end 
          if((cparam_matmul_33_data_stationary == 0) && (matmul_33_row_count >= cparam_matmul_33_max_row_count) && (matmul_33_bat_count >= cparam_matmul_33_max_bat_count) && cparam_matmul_33_keep_input) begin
            matmul_33_skip_read_act <= 1;
          end 
          if((matmul_33_row_count >= cparam_matmul_33_max_row_count) && (matmul_33_bat_count >= cparam_matmul_33_max_bat_count) && (matmul_33_och_count >= cparam_matmul_33_max_och_count)) begin
            matmul_33_skip_comp <= 1;
          end 
          if(matmul_33_skip_write_out && (matmul_33_prev_row_count == 0) && (matmul_33_prev_bat_count == 0) && (matmul_33_prev_och_count == 0)) begin
            matmul_33_skip_write_out <= 0;
          end 
          if(cparam_matmul_33_data_stationary == 0) begin
            control_matmul_33 <= control_matmul_33_12;
          end 
          if((cparam_matmul_33_data_stationary == 0) && (matmul_33_row_count >= cparam_matmul_33_max_row_count) && (matmul_33_bat_count >= cparam_matmul_33_max_bat_count)) begin
            control_matmul_33 <= control_matmul_33_7;
          end 
          if(cparam_matmul_33_data_stationary == 1) begin
            control_matmul_33 <= control_matmul_33_7;
          end 
          if((cparam_matmul_33_data_stationary == 1) && (matmul_33_och_count >= cparam_matmul_33_max_och_count)) begin
            control_matmul_33 <= control_matmul_33_12;
          end 
          if(!matmul_33_skip_write_out && (matmul_33_prev_och_count >= cparam_matmul_33_max_och_count) && (matmul_33_prev_row_count >= cparam_matmul_33_max_row_count) && (matmul_33_prev_bat_count >= cparam_matmul_33_max_bat_count)) begin
            control_matmul_33 <= control_matmul_33_27;
          end 
        end
        control_matmul_33_27: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_matmul_33 <= control_matmul_33_28;
          end 
        end
        control_matmul_33_28: begin
          if(main_fsm == 86) begin
            _control_matmul_33_called <= 0;
          end 
          if(main_fsm == 86) begin
            control_matmul_33 <= control_matmul_33_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_31_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_31 <= write_burst_fsm_31_init;
      write_burst_addr_1636 <= 0;
      write_burst_stride_1637 <= 0;
      write_burst_length_1638 <= 0;
      write_burst_done_1639 <= 0;
    end else begin
      case(write_burst_fsm_31)
        write_burst_fsm_31_init: begin
          write_burst_addr_1636 <= _maxi_read_local_addr_buf;
          write_burst_stride_1637 <= _maxi_read_local_stride_buf;
          write_burst_length_1638 <= _maxi_read_local_size_buf;
          write_burst_done_1639 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 12) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_31 <= write_burst_fsm_31_1;
          end 
        end
        write_burst_fsm_31_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_1636 <= write_burst_addr_1636 + write_burst_stride_1637;
            write_burst_length_1638 <= write_burst_length_1638 - 1;
            write_burst_done_1639 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_1638 <= 1)) begin
            write_burst_done_1639 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_1639 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_1638 <= 1)) begin
            write_burst_fsm_31 <= write_burst_fsm_31_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_31 <= write_burst_fsm_31_init;
          end 
          if(0) begin
            write_burst_fsm_31 <= write_burst_fsm_31_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_32_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_32 <= write_burst_fsm_32_init;
      write_burst_addr_1642 <= 0;
      write_burst_stride_1643 <= 0;
      write_burst_length_1644 <= 0;
      write_burst_done_1645 <= 0;
    end else begin
      case(write_burst_fsm_32)
        write_burst_fsm_32_init: begin
          write_burst_addr_1642 <= _maxi_read_local_addr_buf;
          write_burst_stride_1643 <= _maxi_read_local_stride_buf;
          write_burst_length_1644 <= _maxi_read_local_size_buf;
          write_burst_done_1645 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 13) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_32 <= write_burst_fsm_32_1;
          end 
        end
        write_burst_fsm_32_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_1642 <= write_burst_addr_1642 + write_burst_stride_1643;
            write_burst_length_1644 <= write_burst_length_1644 - 1;
            write_burst_done_1645 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_1644 <= 1)) begin
            write_burst_done_1645 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_1645 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_1644 <= 1)) begin
            write_burst_fsm_32 <= write_burst_fsm_32_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_32 <= write_burst_fsm_32_init;
          end 
          if(0) begin
            write_burst_fsm_32 <= write_burst_fsm_32_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_33_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_33 <= write_burst_fsm_33_init;
      write_burst_addr_1650 <= 0;
      write_burst_stride_1651 <= 0;
      write_burst_length_1652 <= 0;
      write_burst_done_1653 <= 0;
    end else begin
      case(write_burst_fsm_33)
        write_burst_fsm_33_init: begin
          write_burst_addr_1650 <= _maxi_read_local_addr_buf;
          write_burst_stride_1651 <= _maxi_read_local_stride_buf;
          write_burst_length_1652 <= _maxi_read_local_size_buf;
          write_burst_done_1653 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 14) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_33 <= write_burst_fsm_33_1;
          end 
        end
        write_burst_fsm_33_1: begin
          if(write_burst_block_ram_wvalid_1648) begin
            write_burst_addr_1650 <= write_burst_addr_1650 + write_burst_stride_1651;
            write_burst_length_1652 <= write_burst_length_1652 - 1;
            write_burst_done_1653 <= 0;
          end 
          if(write_burst_block_ram_wvalid_1648 && (write_burst_length_1652 <= 1)) begin
            write_burst_done_1653 <= 1;
          end 
          if(write_burst_block_ram_wvalid_1648 && 0) begin
            write_burst_done_1653 <= 1;
          end 
          if(write_burst_block_ram_wvalid_1648 && (write_burst_length_1652 <= 1)) begin
            write_burst_fsm_33 <= write_burst_fsm_33_init;
          end 
          if(write_burst_block_ram_wvalid_1648 && 0) begin
            write_burst_fsm_33 <= write_burst_fsm_33_init;
          end 
          if(write_burst_block_ram_wquit_1649) begin
            write_burst_fsm_33 <= write_burst_fsm_33_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_34_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_34 <= write_burst_fsm_34_init;
      write_burst_addr_1656 <= 0;
      write_burst_stride_1657 <= 0;
      write_burst_length_1658 <= 0;
      write_burst_done_1659 <= 0;
    end else begin
      case(write_burst_fsm_34)
        write_burst_fsm_34_init: begin
          write_burst_addr_1656 <= _maxi_read_local_addr_buf;
          write_burst_stride_1657 <= _maxi_read_local_stride_buf;
          write_burst_length_1658 <= _maxi_read_local_size_buf;
          write_burst_done_1659 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 14) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_34 <= write_burst_fsm_34_1;
          end 
        end
        write_burst_fsm_34_1: begin
          if(write_burst_block_ram_wvalid_1654) begin
            write_burst_addr_1656 <= write_burst_addr_1656 + write_burst_stride_1657;
            write_burst_length_1658 <= write_burst_length_1658 - 1;
            write_burst_done_1659 <= 0;
          end 
          if(write_burst_block_ram_wvalid_1654 && (write_burst_length_1658 <= 1)) begin
            write_burst_done_1659 <= 1;
          end 
          if(write_burst_block_ram_wvalid_1654 && 0) begin
            write_burst_done_1659 <= 1;
          end 
          if(write_burst_block_ram_wvalid_1654 && (write_burst_length_1658 <= 1)) begin
            write_burst_fsm_34 <= write_burst_fsm_34_init;
          end 
          if(write_burst_block_ram_wvalid_1654 && 0) begin
            write_burst_fsm_34 <= write_burst_fsm_34_init;
          end 
          if(write_burst_block_ram_wquit_1655) begin
            write_burst_fsm_34 <= write_burst_fsm_34_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_35_1 = 1;
  localparam write_burst_block_fsm_35_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_35 <= write_burst_block_fsm_35_init;
      write_burst_block_length_1660 <= 0;
      write_burst_block_blocksize_1661 <= 0;
      write_burst_block_done_1662 <= 0;
      write_burst_block_count_1663 <= 0;
    end else begin
      case(write_burst_block_fsm_35)
        write_burst_block_fsm_35_init: begin
          write_burst_block_length_1660 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_1661 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_1662 <= 0;
          write_burst_block_count_1663 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 14) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_35 <= write_burst_block_fsm_35_1;
          end 
        end
        write_burst_block_fsm_35_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_1660 <= write_burst_block_length_1660 - 1;
            write_burst_block_done_1662 <= 0;
            write_burst_block_count_1663 <= write_burst_block_count_1663 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_1660 <= 1)) begin
            write_burst_block_done_1662 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_1662 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_1663 == write_burst_block_blocksize_1661 - 1)) begin
            write_burst_block_count_1663 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_1663 == write_burst_block_blocksize_1661 - 1)) begin
            write_burst_block_fsm_35 <= write_burst_block_fsm_35_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_1660 <= 1)) begin
            write_burst_block_fsm_35 <= write_burst_block_fsm_35_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_35 <= write_burst_block_fsm_35_init;
          end 
          if(0) begin
            write_burst_block_fsm_35 <= write_burst_block_fsm_35_init;
          end 
        end
        write_burst_block_fsm_35_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_1660 <= write_burst_block_length_1660 - 1;
            write_burst_block_done_1662 <= 0;
            write_burst_block_count_1663 <= write_burst_block_count_1663 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_1660 <= 1)) begin
            write_burst_block_done_1662 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_1662 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_1663 == write_burst_block_blocksize_1661 - 1)) begin
            write_burst_block_count_1663 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_1663 == write_burst_block_blocksize_1661 - 1)) begin
            write_burst_block_fsm_35 <= write_burst_block_fsm_35_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_1660 <= 1)) begin
            write_burst_block_fsm_35 <= write_burst_block_fsm_35_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_35 <= write_burst_block_fsm_35_init;
          end 
          if(0) begin
            write_burst_block_fsm_35 <= write_burst_block_fsm_35_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_36_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_36 <= write_burst_fsm_36_init;
      write_burst_addr_1666 <= 0;
      write_burst_stride_1667 <= 0;
      write_burst_length_1668 <= 0;
      write_burst_done_1669 <= 0;
    end else begin
      case(write_burst_fsm_36)
        write_burst_fsm_36_init: begin
          write_burst_addr_1666 <= _maxi_read_local_addr_buf;
          write_burst_stride_1667 <= _maxi_read_local_stride_buf;
          write_burst_length_1668 <= _maxi_read_local_size_buf;
          write_burst_done_1669 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 15) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_36 <= write_burst_fsm_36_1;
          end 
        end
        write_burst_fsm_36_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_1666 <= write_burst_addr_1666 + write_burst_stride_1667;
            write_burst_length_1668 <= write_burst_length_1668 - 1;
            write_burst_done_1669 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_1668 <= 1)) begin
            write_burst_done_1669 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_1669 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_1668 <= 1)) begin
            write_burst_fsm_36 <= write_burst_fsm_36_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_36 <= write_burst_fsm_36_init;
          end 
          if(0) begin
            write_burst_fsm_36 <= write_burst_fsm_36_init;
          end 
        end
      endcase
    end
  end

  localparam matmul_33_comp_fsm_1 = 1;
  localparam matmul_33_comp_fsm_2 = 2;
  localparam matmul_33_comp_fsm_3 = 3;
  localparam matmul_33_comp_fsm_4 = 4;
  localparam matmul_33_comp_fsm_5 = 5;
  localparam matmul_33_comp_fsm_6 = 6;

  always @(posedge CLK) begin
    if(RST) begin
      matmul_33_comp_fsm <= matmul_33_comp_fsm_init;
      matmul_33_stream_act_local_0 <= 0;
      matmul_33_stream_out_local_col <= 0;
      matmul_33_stream_out_local_val <= 0;
      matmul_33_col_count <= 0;
      matmul_33_col_select <= 0;
      matmul_33_filter_page_comp_offset_buf <= 0;
      matmul_33_act_page_comp_offset_buf_0 <= 0;
      matmul_33_out_page_comp_offset_buf <= 0;
      matmul_33_row_count_buf <= 0;
      matmul_33_row_select_buf <= 0;
      matmul_33_och_count_buf <= 0;
      matmul_33_next_stream_num_ops <= 0;
      matmul_33_stream_pad_masks <= 0;
      matmul_33_sync_comp_count <= 0;
    end else begin
      if(_stream_matmul_33_sink_stop) begin
        matmul_33_sync_comp_count <= matmul_33_sync_comp_count + 1;
      end 
      if(control_matmul_33 == 6) begin
        matmul_33_sync_comp_count <= 0;
      end 
      case(matmul_33_comp_fsm)
        matmul_33_comp_fsm_init: begin
          if((control_matmul_33 == 19) && !matmul_33_skip_comp) begin
            matmul_33_comp_fsm <= matmul_33_comp_fsm_1;
          end 
        end
        matmul_33_comp_fsm_1: begin
          matmul_33_stream_act_local_0 <= 0;
          if(cparam_matmul_33_stream_act_local_small_flags_0) begin
            matmul_33_stream_act_local_0 <= cparam_matmul_33_stream_act_local_small_offset;
          end 
          if(cparam_matmul_33_stream_act_local_large_flags_0) begin
            matmul_33_stream_act_local_0 <= cparam_matmul_33_stream_act_local_large_offset;
          end 
          matmul_33_stream_out_local_col <= 0;
          if((cparam_matmul_33_data_stationary == 1) && (matmul_33_och_count == 0)) begin
            matmul_33_stream_out_local_val <= 0;
          end 
          matmul_33_col_count <= 0;
          matmul_33_col_select <= cparam_matmul_33_col_select_initval;
          matmul_33_filter_page_comp_offset_buf <= matmul_33_filter_page_comp_offset;
          matmul_33_act_page_comp_offset_buf_0 <= matmul_33_act_page_comp_offset_0;
          matmul_33_out_page_comp_offset_buf <= matmul_33_out_page_comp_offset;
          matmul_33_row_count_buf <= matmul_33_row_count;
          matmul_33_row_select_buf <= matmul_33_row_select;
          matmul_33_och_count_buf <= matmul_33_och_count;
          matmul_33_next_stream_num_ops <= (matmul_33_och_count >= cparam_matmul_33_max_och_count)? cparam_matmul_33_stream_num_ops_res : cparam_matmul_33_stream_num_ops;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_2;
        end
        matmul_33_comp_fsm_2: begin
          matmul_33_stream_pad_masks <= { matmul_33_stream_pad_mask_0_0 };
          matmul_33_comp_fsm <= matmul_33_comp_fsm_3;
        end
        matmul_33_comp_fsm_3: begin
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          if(_stream_matmul_33_stream_oready) begin
            matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
          end 
          matmul_33_comp_fsm <= matmul_33_comp_fsm_4;
        end
        matmul_33_comp_fsm_4: begin
          if(!_stream_matmul_33_source_busy) begin
            matmul_33_comp_fsm <= matmul_33_comp_fsm_5;
          end 
        end
        matmul_33_comp_fsm_5: begin
          if(_stream_matmul_33_busy) begin
            matmul_33_comp_fsm <= matmul_33_comp_fsm_6;
          end 
        end
        matmul_33_comp_fsm_6: begin
          if(!((matmul_33_col_select == 0)? cparam_matmul_33_inc_act_laddr_conds_0 : 0)) begin
            matmul_33_stream_act_local_0 <= matmul_33_stream_act_local_0 + cparam_matmul_33_inc_act_laddr_small;
          end 
          if((matmul_33_col_select == 0)? cparam_matmul_33_inc_act_laddr_conds_0 : 0) begin
            matmul_33_stream_act_local_0 <= matmul_33_stream_act_local_0 + cparam_matmul_33_inc_act_laddr_large;
          end 
          if(matmul_33_col_count >= cparam_matmul_33_max_col_count) begin
            matmul_33_stream_act_local_0 <= 0;
          end 
          if((matmul_33_col_count >= cparam_matmul_33_max_col_count) && cparam_matmul_33_stream_act_local_small_flags_0) begin
            matmul_33_stream_act_local_0 <= cparam_matmul_33_stream_act_local_small_offset;
          end 
          if((matmul_33_col_count >= cparam_matmul_33_max_col_count) && cparam_matmul_33_stream_act_local_large_flags_0) begin
            matmul_33_stream_act_local_0 <= cparam_matmul_33_stream_act_local_large_offset;
          end 
          if(cparam_matmul_33_data_stationary == 0) begin
            matmul_33_stream_out_local_col <= matmul_33_stream_out_local_col + matmul_33_next_stream_num_ops;
          end 
          if((cparam_matmul_33_data_stationary == 0) && (matmul_33_col_count >= cparam_matmul_33_max_col_count)) begin
            matmul_33_stream_out_local_col <= 0;
          end 
          if(cparam_matmul_33_data_stationary == 1) begin
            matmul_33_stream_out_local_col <= matmul_33_stream_out_local_col + cparam_matmul_33_inc_out_laddr_col;
          end 
          if((cparam_matmul_33_data_stationary == 1) && (matmul_33_col_count >= cparam_matmul_33_max_col_count)) begin
            matmul_33_stream_out_local_val <= matmul_33_stream_out_local_val + matmul_33_next_stream_num_ops;
            matmul_33_stream_out_local_col <= 0;
          end 
          matmul_33_col_count <= matmul_33_col_count + cparam_matmul_33_stride_col_par_col;
          if(matmul_33_col_count >= cparam_matmul_33_max_col_count) begin
            matmul_33_col_count <= 0;
          end 
          matmul_33_col_select <= matmul_33_col_select + cparam_matmul_33_stride_col_mod_filter_num;
          if(matmul_33_col_select + cparam_matmul_33_stride_col_mod_filter_num >= 1) begin
            matmul_33_col_select <= matmul_33_col_select - cparam_matmul_33_filter_num_col_minus_stride_col_mod;
          end 
          if(matmul_33_col_count >= cparam_matmul_33_max_col_count) begin
            matmul_33_col_select <= cparam_matmul_33_col_select_initval;
          end 
          matmul_33_comp_fsm <= matmul_33_comp_fsm_2;
          if(matmul_33_col_count >= cparam_matmul_33_max_col_count) begin
            matmul_33_comp_fsm <= matmul_33_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_33_source_7_source_pat_fsm_0_1 = 1;
  localparam _stream_matmul_33_source_7_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_33_source_7_source_pat_fsm_0 <= _stream_matmul_33_source_7_source_pat_fsm_0_init;
    end else begin
      case(_stream_matmul_33_source_7_source_pat_fsm_0)
        _stream_matmul_33_source_7_source_pat_fsm_0_init: begin
          if(_stream_matmul_33_source_start && _stream_matmul_33_source_7_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_7_source_pat_fsm_0 <= _stream_matmul_33_source_7_source_pat_fsm_0_1;
          end 
        end
        _stream_matmul_33_source_7_source_pat_fsm_0_1: begin
          if(_stream_matmul_33_source_stop && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_7_source_pat_fsm_0 <= _stream_matmul_33_source_7_source_pat_fsm_0_init;
          end 
          if((_source_stream_matmul_33_source_7_pat_count_0 == 0) && (_source_stream_matmul_33_source_7_pat_count_1 == 0) && (_source_stream_matmul_33_source_7_pat_count_2 == 0) && (_source_stream_matmul_33_source_7_pat_count_3 == 0) && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_7_source_pat_fsm_0 <= _stream_matmul_33_source_7_source_pat_fsm_0_2;
          end 
        end
        _stream_matmul_33_source_7_source_pat_fsm_0_2: begin
          if(_stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_7_source_pat_fsm_0 <= _stream_matmul_33_source_7_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_33_source_9_source_pat_fsm_1_1 = 1;
  localparam _stream_matmul_33_source_9_source_pat_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_33_source_9_source_pat_fsm_1 <= _stream_matmul_33_source_9_source_pat_fsm_1_init;
    end else begin
      case(_stream_matmul_33_source_9_source_pat_fsm_1)
        _stream_matmul_33_source_9_source_pat_fsm_1_init: begin
          if(_stream_matmul_33_source_start && _stream_matmul_33_source_9_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_9_source_pat_fsm_1 <= _stream_matmul_33_source_9_source_pat_fsm_1_1;
          end 
        end
        _stream_matmul_33_source_9_source_pat_fsm_1_1: begin
          if(_stream_matmul_33_source_stop && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_9_source_pat_fsm_1 <= _stream_matmul_33_source_9_source_pat_fsm_1_init;
          end 
          if((_source_stream_matmul_33_source_9_pat_count_0 == 0) && (_source_stream_matmul_33_source_9_pat_count_1 == 0) && (_source_stream_matmul_33_source_9_pat_count_2 == 0) && (_source_stream_matmul_33_source_9_pat_count_3 == 0) && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_9_source_pat_fsm_1 <= _stream_matmul_33_source_9_source_pat_fsm_1_2;
          end 
        end
        _stream_matmul_33_source_9_source_pat_fsm_1_2: begin
          if(_stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_9_source_pat_fsm_1 <= _stream_matmul_33_source_9_source_pat_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_33_source_20_source_pat_fsm_2_1 = 1;
  localparam _stream_matmul_33_source_20_source_pat_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_33_source_20_source_pat_fsm_2 <= _stream_matmul_33_source_20_source_pat_fsm_2_init;
    end else begin
      case(_stream_matmul_33_source_20_source_pat_fsm_2)
        _stream_matmul_33_source_20_source_pat_fsm_2_init: begin
          if(_stream_matmul_33_source_start && _stream_matmul_33_source_20_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_20_source_pat_fsm_2 <= _stream_matmul_33_source_20_source_pat_fsm_2_1;
          end 
        end
        _stream_matmul_33_source_20_source_pat_fsm_2_1: begin
          if(_stream_matmul_33_source_stop && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_20_source_pat_fsm_2 <= _stream_matmul_33_source_20_source_pat_fsm_2_init;
          end 
          if((_source_stream_matmul_33_source_20_pat_count_0 == 0) && (_source_stream_matmul_33_source_20_pat_count_1 == 0) && (_source_stream_matmul_33_source_20_pat_count_2 == 0) && (_source_stream_matmul_33_source_20_pat_count_3 == 0) && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_20_source_pat_fsm_2 <= _stream_matmul_33_source_20_source_pat_fsm_2_2;
          end 
        end
        _stream_matmul_33_source_20_source_pat_fsm_2_2: begin
          if(_stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_20_source_pat_fsm_2 <= _stream_matmul_33_source_20_source_pat_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_33_source_21_source_pat_fsm_3_1 = 1;
  localparam _stream_matmul_33_source_21_source_pat_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_33_source_21_source_pat_fsm_3 <= _stream_matmul_33_source_21_source_pat_fsm_3_init;
    end else begin
      case(_stream_matmul_33_source_21_source_pat_fsm_3)
        _stream_matmul_33_source_21_source_pat_fsm_3_init: begin
          if(_stream_matmul_33_source_start && _stream_matmul_33_source_21_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_21_source_pat_fsm_3 <= _stream_matmul_33_source_21_source_pat_fsm_3_1;
          end 
        end
        _stream_matmul_33_source_21_source_pat_fsm_3_1: begin
          if(_stream_matmul_33_source_stop && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_21_source_pat_fsm_3 <= _stream_matmul_33_source_21_source_pat_fsm_3_init;
          end 
          if((_source_stream_matmul_33_source_21_pat_count_0 == 0) && (_source_stream_matmul_33_source_21_pat_count_1 == 0) && (_source_stream_matmul_33_source_21_pat_count_2 == 0) && (_source_stream_matmul_33_source_21_pat_count_3 == 0) && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_21_source_pat_fsm_3 <= _stream_matmul_33_source_21_source_pat_fsm_3_2;
          end 
        end
        _stream_matmul_33_source_21_source_pat_fsm_3_2: begin
          if(_stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_21_source_pat_fsm_3 <= _stream_matmul_33_source_21_source_pat_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_33_source_22_source_pat_fsm_4_1 = 1;
  localparam _stream_matmul_33_source_22_source_pat_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_33_source_22_source_pat_fsm_4 <= _stream_matmul_33_source_22_source_pat_fsm_4_init;
    end else begin
      case(_stream_matmul_33_source_22_source_pat_fsm_4)
        _stream_matmul_33_source_22_source_pat_fsm_4_init: begin
          if(_stream_matmul_33_source_start && _stream_matmul_33_source_22_source_mode & 5'b10 && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_22_source_pat_fsm_4 <= _stream_matmul_33_source_22_source_pat_fsm_4_1;
          end 
        end
        _stream_matmul_33_source_22_source_pat_fsm_4_1: begin
          if(_stream_matmul_33_source_stop && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_22_source_pat_fsm_4 <= _stream_matmul_33_source_22_source_pat_fsm_4_init;
          end 
          if((_source_stream_matmul_33_source_22_pat_count_0 == 0) && (_source_stream_matmul_33_source_22_pat_count_1 == 0) && (_source_stream_matmul_33_source_22_pat_count_2 == 0) && (_source_stream_matmul_33_source_22_pat_count_3 == 0) && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_22_source_pat_fsm_4 <= _stream_matmul_33_source_22_source_pat_fsm_4_2;
          end 
        end
        _stream_matmul_33_source_22_source_pat_fsm_4_2: begin
          if(_stream_matmul_33_stream_oready) begin
            _stream_matmul_33_source_22_source_pat_fsm_4 <= _stream_matmul_33_source_22_source_pat_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_33_sink_33_sink_fsm_5_1 = 1;
  localparam _stream_matmul_33_sink_33_sink_fsm_5_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_33_sink_33_sink_fsm_5 <= _stream_matmul_33_sink_33_sink_fsm_5_init;
    end else begin
      case(_stream_matmul_33_sink_33_sink_fsm_5)
        _stream_matmul_33_sink_33_sink_fsm_5_init: begin
          if(_stream_matmul_33_sink_start && _stream_matmul_33_sink_33_sink_mode & 5'b1 && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_sink_33_sink_fsm_5 <= _stream_matmul_33_sink_33_sink_fsm_5_1;
          end 
        end
        _stream_matmul_33_sink_33_sink_fsm_5_1: begin
          if(_stream_matmul_33_stream_oready) begin
            _stream_matmul_33_sink_33_sink_fsm_5 <= _stream_matmul_33_sink_33_sink_fsm_5_2;
          end 
        end
        _stream_matmul_33_sink_33_sink_fsm_5_2: begin
          if(stream_matmul_33_sink_34_data && (_stream_matmul_33_sink_33_sink_count == 1) && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_sink_33_sink_fsm_5 <= _stream_matmul_33_sink_33_sink_fsm_5_init;
          end 
          if(_stream_matmul_33_sink_stop && _stream_matmul_33_stream_oready) begin
            _stream_matmul_33_sink_33_sink_fsm_5 <= _stream_matmul_33_sink_33_sink_fsm_5_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_fsm_37_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_fsm_37 <= read_burst_fsm_37_init;
      read_burst_addr_2009 <= 0;
      read_burst_stride_2010 <= 0;
      read_burst_length_2011 <= 0;
      read_burst_rvalid_2012 <= 0;
      read_burst_rlast_2013 <= 0;
    end else begin
      case(read_burst_fsm_37)
        read_burst_fsm_37_init: begin
          read_burst_addr_2009 <= _maxi_write_local_addr_buf;
          read_burst_stride_2010 <= _maxi_write_local_stride_buf;
          read_burst_length_2011 <= _maxi_write_size_buf;
          read_burst_rvalid_2012 <= 0;
          read_burst_rlast_2013 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 3) && (_maxi_write_size_buf > 0)) begin
            read_burst_fsm_37 <= read_burst_fsm_37_1;
          end 
        end
        read_burst_fsm_37_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_2011 > 0)) begin
            read_burst_addr_2009 <= read_burst_addr_2009 + read_burst_stride_2010;
            read_burst_length_2011 <= read_burst_length_2011 - 1;
            read_burst_rvalid_2012 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_2011 <= 1)) begin
            read_burst_rlast_2013 <= 1;
          end 
          if(read_burst_rlast_2013 && read_burst_rvalid_2012 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_rvalid_2012 <= 0;
            read_burst_rlast_2013 <= 0;
          end 
          if(0) begin
            read_burst_rvalid_2012 <= 0;
            read_burst_rlast_2013 <= 0;
          end 
          if(read_burst_rlast_2013 && read_burst_rvalid_2012 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_fsm_37 <= read_burst_fsm_37_init;
          end 
          if(0) begin
            read_burst_fsm_37 <= read_burst_fsm_37_init;
          end 
        end
      endcase
    end
  end


endmodule



module _maxi_read_req_fifo
(
  input CLK,
  input RST,
  input _maxi_read_req_fifo_enq,
  input [137-1:0] _maxi_read_req_fifo_wdata,
  output _maxi_read_req_fifo_full,
  output _maxi_read_req_fifo_almost_full,
  input _maxi_read_req_fifo_deq,
  output [137-1:0] _maxi_read_req_fifo_rdata,
  output _maxi_read_req_fifo_empty,
  output _maxi_read_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _maxi_read_req_fifo_full = is_full;
  assign _maxi_read_req_fifo_almost_full = is_almost_full || is_full;
  assign _maxi_read_req_fifo_empty = is_empty;
  assign _maxi_read_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _maxi_read_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_maxi_read_req_fifo_enq && !is_full) begin
        mem[head] <= _maxi_read_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_maxi_read_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module _maxi_write_req_fifo
(
  input CLK,
  input RST,
  input _maxi_write_req_fifo_enq,
  input [137-1:0] _maxi_write_req_fifo_wdata,
  output _maxi_write_req_fifo_full,
  output _maxi_write_req_fifo_almost_full,
  input _maxi_write_req_fifo_deq,
  output [137-1:0] _maxi_write_req_fifo_rdata,
  output _maxi_write_req_fifo_empty,
  output _maxi_write_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _maxi_write_req_fifo_full = is_full;
  assign _maxi_write_req_fifo_almost_full = is_almost_full || is_full;
  assign _maxi_write_req_fifo_empty = is_empty;
  assign _maxi_write_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _maxi_write_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_maxi_write_req_fifo_enq && !is_full) begin
        mem[head] <= _maxi_write_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_maxi_write_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module ram_w16_l16384_id0_0
(
  input CLK,
  input [13-1:0] ram_w16_l16384_id0_0_0_addr,
  output [16-1:0] ram_w16_l16384_id0_0_0_rdata,
  input [16-1:0] ram_w16_l16384_id0_0_0_wdata,
  input ram_w16_l16384_id0_0_0_wenable,
  input ram_w16_l16384_id0_0_0_enable,
  input [13-1:0] ram_w16_l16384_id0_0_1_addr,
  output [16-1:0] ram_w16_l16384_id0_0_1_rdata,
  input [16-1:0] ram_w16_l16384_id0_0_1_wdata,
  input ram_w16_l16384_id0_0_1_wenable,
  input ram_w16_l16384_id0_0_1_enable
);

  reg [16-1:0] ram_w16_l16384_id0_0_0_rdata_out;
  assign ram_w16_l16384_id0_0_0_rdata = ram_w16_l16384_id0_0_0_rdata_out;
  reg [16-1:0] ram_w16_l16384_id0_0_1_rdata_out;
  assign ram_w16_l16384_id0_0_1_rdata = ram_w16_l16384_id0_0_1_rdata_out;
  reg [16-1:0] mem [0:8192-1];

  always @(posedge CLK) begin
    if(ram_w16_l16384_id0_0_0_enable) begin
      if(ram_w16_l16384_id0_0_0_wenable) begin
        mem[ram_w16_l16384_id0_0_0_addr] <= ram_w16_l16384_id0_0_0_wdata;
        ram_w16_l16384_id0_0_0_rdata_out <= ram_w16_l16384_id0_0_0_wdata;
      end else begin
        ram_w16_l16384_id0_0_0_rdata_out <= mem[ram_w16_l16384_id0_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l16384_id0_0_1_enable) begin
      if(ram_w16_l16384_id0_0_1_wenable) begin
        mem[ram_w16_l16384_id0_0_1_addr] <= ram_w16_l16384_id0_0_1_wdata;
        ram_w16_l16384_id0_0_1_rdata_out <= ram_w16_l16384_id0_0_1_wdata;
      end else begin
        ram_w16_l16384_id0_0_1_rdata_out <= mem[ram_w16_l16384_id0_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l16384_id0_1
(
  input CLK,
  input [13-1:0] ram_w16_l16384_id0_1_0_addr,
  output [16-1:0] ram_w16_l16384_id0_1_0_rdata,
  input [16-1:0] ram_w16_l16384_id0_1_0_wdata,
  input ram_w16_l16384_id0_1_0_wenable,
  input ram_w16_l16384_id0_1_0_enable,
  input [13-1:0] ram_w16_l16384_id0_1_1_addr,
  output [16-1:0] ram_w16_l16384_id0_1_1_rdata,
  input [16-1:0] ram_w16_l16384_id0_1_1_wdata,
  input ram_w16_l16384_id0_1_1_wenable,
  input ram_w16_l16384_id0_1_1_enable
);

  reg [16-1:0] ram_w16_l16384_id0_1_0_rdata_out;
  assign ram_w16_l16384_id0_1_0_rdata = ram_w16_l16384_id0_1_0_rdata_out;
  reg [16-1:0] ram_w16_l16384_id0_1_1_rdata_out;
  assign ram_w16_l16384_id0_1_1_rdata = ram_w16_l16384_id0_1_1_rdata_out;
  reg [16-1:0] mem [0:8192-1];

  always @(posedge CLK) begin
    if(ram_w16_l16384_id0_1_0_enable) begin
      if(ram_w16_l16384_id0_1_0_wenable) begin
        mem[ram_w16_l16384_id0_1_0_addr] <= ram_w16_l16384_id0_1_0_wdata;
        ram_w16_l16384_id0_1_0_rdata_out <= ram_w16_l16384_id0_1_0_wdata;
      end else begin
        ram_w16_l16384_id0_1_0_rdata_out <= mem[ram_w16_l16384_id0_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l16384_id0_1_1_enable) begin
      if(ram_w16_l16384_id0_1_1_wenable) begin
        mem[ram_w16_l16384_id0_1_1_addr] <= ram_w16_l16384_id0_1_1_wdata;
        ram_w16_l16384_id0_1_1_rdata_out <= ram_w16_l16384_id0_1_1_wdata;
      end else begin
        ram_w16_l16384_id0_1_1_rdata_out <= mem[ram_w16_l16384_id0_1_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l4096_id0
(
  input CLK,
  input [12-1:0] ram_w32_l4096_id0_0_addr,
  output [32-1:0] ram_w32_l4096_id0_0_rdata,
  input [32-1:0] ram_w32_l4096_id0_0_wdata,
  input ram_w32_l4096_id0_0_wenable,
  input ram_w32_l4096_id0_0_enable,
  input [12-1:0] ram_w32_l4096_id0_1_addr,
  output [32-1:0] ram_w32_l4096_id0_1_rdata,
  input [32-1:0] ram_w32_l4096_id0_1_wdata,
  input ram_w32_l4096_id0_1_wenable,
  input ram_w32_l4096_id0_1_enable
);

  reg [32-1:0] ram_w32_l4096_id0_0_rdata_out;
  assign ram_w32_l4096_id0_0_rdata = ram_w32_l4096_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l4096_id0_1_rdata_out;
  assign ram_w32_l4096_id0_1_rdata = ram_w32_l4096_id0_1_rdata_out;
  reg [32-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w32_l4096_id0_0_enable) begin
      if(ram_w32_l4096_id0_0_wenable) begin
        mem[ram_w32_l4096_id0_0_addr] <= ram_w32_l4096_id0_0_wdata;
        ram_w32_l4096_id0_0_rdata_out <= ram_w32_l4096_id0_0_wdata;
      end else begin
        ram_w32_l4096_id0_0_rdata_out <= mem[ram_w32_l4096_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l4096_id0_1_enable) begin
      if(ram_w32_l4096_id0_1_wenable) begin
        mem[ram_w32_l4096_id0_1_addr] <= ram_w32_l4096_id0_1_wdata;
        ram_w32_l4096_id0_1_rdata_out <= ram_w32_l4096_id0_1_wdata;
      end else begin
        ram_w32_l4096_id0_1_rdata_out <= mem[ram_w32_l4096_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l4096_id0_0
(
  input CLK,
  input [11-1:0] ram_w16_l4096_id0_0_0_addr,
  output [16-1:0] ram_w16_l4096_id0_0_0_rdata,
  input [16-1:0] ram_w16_l4096_id0_0_0_wdata,
  input ram_w16_l4096_id0_0_0_wenable,
  input ram_w16_l4096_id0_0_0_enable,
  input [11-1:0] ram_w16_l4096_id0_0_1_addr,
  output [16-1:0] ram_w16_l4096_id0_0_1_rdata,
  input [16-1:0] ram_w16_l4096_id0_0_1_wdata,
  input ram_w16_l4096_id0_0_1_wenable,
  input ram_w16_l4096_id0_0_1_enable
);

  reg [16-1:0] ram_w16_l4096_id0_0_0_rdata_out;
  assign ram_w16_l4096_id0_0_0_rdata = ram_w16_l4096_id0_0_0_rdata_out;
  reg [16-1:0] ram_w16_l4096_id0_0_1_rdata_out;
  assign ram_w16_l4096_id0_0_1_rdata = ram_w16_l4096_id0_0_1_rdata_out;
  reg [16-1:0] mem [0:2048-1];

  always @(posedge CLK) begin
    if(ram_w16_l4096_id0_0_0_enable) begin
      if(ram_w16_l4096_id0_0_0_wenable) begin
        mem[ram_w16_l4096_id0_0_0_addr] <= ram_w16_l4096_id0_0_0_wdata;
        ram_w16_l4096_id0_0_0_rdata_out <= ram_w16_l4096_id0_0_0_wdata;
      end else begin
        ram_w16_l4096_id0_0_0_rdata_out <= mem[ram_w16_l4096_id0_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l4096_id0_0_1_enable) begin
      if(ram_w16_l4096_id0_0_1_wenable) begin
        mem[ram_w16_l4096_id0_0_1_addr] <= ram_w16_l4096_id0_0_1_wdata;
        ram_w16_l4096_id0_0_1_rdata_out <= ram_w16_l4096_id0_0_1_wdata;
      end else begin
        ram_w16_l4096_id0_0_1_rdata_out <= mem[ram_w16_l4096_id0_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l4096_id0_1
(
  input CLK,
  input [11-1:0] ram_w16_l4096_id0_1_0_addr,
  output [16-1:0] ram_w16_l4096_id0_1_0_rdata,
  input [16-1:0] ram_w16_l4096_id0_1_0_wdata,
  input ram_w16_l4096_id0_1_0_wenable,
  input ram_w16_l4096_id0_1_0_enable,
  input [11-1:0] ram_w16_l4096_id0_1_1_addr,
  output [16-1:0] ram_w16_l4096_id0_1_1_rdata,
  input [16-1:0] ram_w16_l4096_id0_1_1_wdata,
  input ram_w16_l4096_id0_1_1_wenable,
  input ram_w16_l4096_id0_1_1_enable
);

  reg [16-1:0] ram_w16_l4096_id0_1_0_rdata_out;
  assign ram_w16_l4096_id0_1_0_rdata = ram_w16_l4096_id0_1_0_rdata_out;
  reg [16-1:0] ram_w16_l4096_id0_1_1_rdata_out;
  assign ram_w16_l4096_id0_1_1_rdata = ram_w16_l4096_id0_1_1_rdata_out;
  reg [16-1:0] mem [0:2048-1];

  always @(posedge CLK) begin
    if(ram_w16_l4096_id0_1_0_enable) begin
      if(ram_w16_l4096_id0_1_0_wenable) begin
        mem[ram_w16_l4096_id0_1_0_addr] <= ram_w16_l4096_id0_1_0_wdata;
        ram_w16_l4096_id0_1_0_rdata_out <= ram_w16_l4096_id0_1_0_wdata;
      end else begin
        ram_w16_l4096_id0_1_0_rdata_out <= mem[ram_w16_l4096_id0_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l4096_id0_1_1_enable) begin
      if(ram_w16_l4096_id0_1_1_wenable) begin
        mem[ram_w16_l4096_id0_1_1_addr] <= ram_w16_l4096_id0_1_1_wdata;
        ram_w16_l4096_id0_1_1_rdata_out <= ram_w16_l4096_id0_1_1_wdata;
      end else begin
        ram_w16_l4096_id0_1_1_rdata_out <= mem[ram_w16_l4096_id0_1_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l1024_id0
(
  input CLK,
  input [10-1:0] ram_w32_l1024_id0_0_addr,
  output [32-1:0] ram_w32_l1024_id0_0_rdata,
  input [32-1:0] ram_w32_l1024_id0_0_wdata,
  input ram_w32_l1024_id0_0_wenable,
  input ram_w32_l1024_id0_0_enable,
  input [10-1:0] ram_w32_l1024_id0_1_addr,
  output [32-1:0] ram_w32_l1024_id0_1_rdata,
  input [32-1:0] ram_w32_l1024_id0_1_wdata,
  input ram_w32_l1024_id0_1_wenable,
  input ram_w32_l1024_id0_1_enable
);

  reg [32-1:0] ram_w32_l1024_id0_0_rdata_out;
  assign ram_w32_l1024_id0_0_rdata = ram_w32_l1024_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l1024_id0_1_rdata_out;
  assign ram_w32_l1024_id0_1_rdata = ram_w32_l1024_id0_1_rdata_out;
  reg [32-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w32_l1024_id0_0_enable) begin
      if(ram_w32_l1024_id0_0_wenable) begin
        mem[ram_w32_l1024_id0_0_addr] <= ram_w32_l1024_id0_0_wdata;
        ram_w32_l1024_id0_0_rdata_out <= ram_w32_l1024_id0_0_wdata;
      end else begin
        ram_w32_l1024_id0_0_rdata_out <= mem[ram_w32_l1024_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l1024_id0_1_enable) begin
      if(ram_w32_l1024_id0_1_wenable) begin
        mem[ram_w32_l1024_id0_1_addr] <= ram_w32_l1024_id0_1_wdata;
        ram_w32_l1024_id0_1_rdata_out <= ram_w32_l1024_id0_1_wdata;
      end else begin
        ram_w32_l1024_id0_1_rdata_out <= mem[ram_w32_l1024_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l512_id0
(
  input CLK,
  input [9-1:0] ram_w32_l512_id0_0_addr,
  output [32-1:0] ram_w32_l512_id0_0_rdata,
  input [32-1:0] ram_w32_l512_id0_0_wdata,
  input ram_w32_l512_id0_0_wenable,
  input ram_w32_l512_id0_0_enable,
  input [9-1:0] ram_w32_l512_id0_1_addr,
  output [32-1:0] ram_w32_l512_id0_1_rdata,
  input [32-1:0] ram_w32_l512_id0_1_wdata,
  input ram_w32_l512_id0_1_wenable,
  input ram_w32_l512_id0_1_enable
);

  reg [32-1:0] ram_w32_l512_id0_0_rdata_out;
  assign ram_w32_l512_id0_0_rdata = ram_w32_l512_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l512_id0_1_rdata_out;
  assign ram_w32_l512_id0_1_rdata = ram_w32_l512_id0_1_rdata_out;
  reg [32-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w32_l512_id0_0_enable) begin
      if(ram_w32_l512_id0_0_wenable) begin
        mem[ram_w32_l512_id0_0_addr] <= ram_w32_l512_id0_0_wdata;
        ram_w32_l512_id0_0_rdata_out <= ram_w32_l512_id0_0_wdata;
      end else begin
        ram_w32_l512_id0_0_rdata_out <= mem[ram_w32_l512_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l512_id0_1_enable) begin
      if(ram_w32_l512_id0_1_wenable) begin
        mem[ram_w32_l512_id0_1_addr] <= ram_w32_l512_id0_1_wdata;
        ram_w32_l512_id0_1_rdata_out <= ram_w32_l512_id0_1_wdata;
      end else begin
        ram_w32_l512_id0_1_rdata_out <= mem[ram_w32_l512_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l512_id1
(
  input CLK,
  input [9-1:0] ram_w32_l512_id1_0_addr,
  output [32-1:0] ram_w32_l512_id1_0_rdata,
  input [32-1:0] ram_w32_l512_id1_0_wdata,
  input ram_w32_l512_id1_0_wenable,
  input ram_w32_l512_id1_0_enable,
  input [9-1:0] ram_w32_l512_id1_1_addr,
  output [32-1:0] ram_w32_l512_id1_1_rdata,
  input [32-1:0] ram_w32_l512_id1_1_wdata,
  input ram_w32_l512_id1_1_wenable,
  input ram_w32_l512_id1_1_enable
);

  reg [32-1:0] ram_w32_l512_id1_0_rdata_out;
  assign ram_w32_l512_id1_0_rdata = ram_w32_l512_id1_0_rdata_out;
  reg [32-1:0] ram_w32_l512_id1_1_rdata_out;
  assign ram_w32_l512_id1_1_rdata = ram_w32_l512_id1_1_rdata_out;
  reg [32-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w32_l512_id1_0_enable) begin
      if(ram_w32_l512_id1_0_wenable) begin
        mem[ram_w32_l512_id1_0_addr] <= ram_w32_l512_id1_0_wdata;
        ram_w32_l512_id1_0_rdata_out <= ram_w32_l512_id1_0_wdata;
      end else begin
        ram_w32_l512_id1_0_rdata_out <= mem[ram_w32_l512_id1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l512_id1_1_enable) begin
      if(ram_w32_l512_id1_1_wenable) begin
        mem[ram_w32_l512_id1_1_addr] <= ram_w32_l512_id1_1_wdata;
        ram_w32_l512_id1_1_rdata_out <= ram_w32_l512_id1_1_wdata;
      end else begin
        ram_w32_l512_id1_1_rdata_out <= mem[ram_w32_l512_id1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id0_0
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id0_0_0_addr,
  output [16-1:0] ram_w16_l1024_id0_0_0_rdata,
  input [16-1:0] ram_w16_l1024_id0_0_0_wdata,
  input ram_w16_l1024_id0_0_0_wenable,
  input ram_w16_l1024_id0_0_0_enable,
  input [9-1:0] ram_w16_l1024_id0_0_1_addr,
  output [16-1:0] ram_w16_l1024_id0_0_1_rdata,
  input [16-1:0] ram_w16_l1024_id0_0_1_wdata,
  input ram_w16_l1024_id0_0_1_wenable,
  input ram_w16_l1024_id0_0_1_enable
);

  reg [16-1:0] ram_w16_l1024_id0_0_0_rdata_out;
  assign ram_w16_l1024_id0_0_0_rdata = ram_w16_l1024_id0_0_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id0_0_1_rdata_out;
  assign ram_w16_l1024_id0_0_1_rdata = ram_w16_l1024_id0_0_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id0_0_0_enable) begin
      if(ram_w16_l1024_id0_0_0_wenable) begin
        mem[ram_w16_l1024_id0_0_0_addr] <= ram_w16_l1024_id0_0_0_wdata;
        ram_w16_l1024_id0_0_0_rdata_out <= ram_w16_l1024_id0_0_0_wdata;
      end else begin
        ram_w16_l1024_id0_0_0_rdata_out <= mem[ram_w16_l1024_id0_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id0_0_1_enable) begin
      if(ram_w16_l1024_id0_0_1_wenable) begin
        mem[ram_w16_l1024_id0_0_1_addr] <= ram_w16_l1024_id0_0_1_wdata;
        ram_w16_l1024_id0_0_1_rdata_out <= ram_w16_l1024_id0_0_1_wdata;
      end else begin
        ram_w16_l1024_id0_0_1_rdata_out <= mem[ram_w16_l1024_id0_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id0_1
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id0_1_0_addr,
  output [16-1:0] ram_w16_l1024_id0_1_0_rdata,
  input [16-1:0] ram_w16_l1024_id0_1_0_wdata,
  input ram_w16_l1024_id0_1_0_wenable,
  input ram_w16_l1024_id0_1_0_enable,
  input [9-1:0] ram_w16_l1024_id0_1_1_addr,
  output [16-1:0] ram_w16_l1024_id0_1_1_rdata,
  input [16-1:0] ram_w16_l1024_id0_1_1_wdata,
  input ram_w16_l1024_id0_1_1_wenable,
  input ram_w16_l1024_id0_1_1_enable
);

  reg [16-1:0] ram_w16_l1024_id0_1_0_rdata_out;
  assign ram_w16_l1024_id0_1_0_rdata = ram_w16_l1024_id0_1_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id0_1_1_rdata_out;
  assign ram_w16_l1024_id0_1_1_rdata = ram_w16_l1024_id0_1_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id0_1_0_enable) begin
      if(ram_w16_l1024_id0_1_0_wenable) begin
        mem[ram_w16_l1024_id0_1_0_addr] <= ram_w16_l1024_id0_1_0_wdata;
        ram_w16_l1024_id0_1_0_rdata_out <= ram_w16_l1024_id0_1_0_wdata;
      end else begin
        ram_w16_l1024_id0_1_0_rdata_out <= mem[ram_w16_l1024_id0_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id0_1_1_enable) begin
      if(ram_w16_l1024_id0_1_1_wenable) begin
        mem[ram_w16_l1024_id0_1_1_addr] <= ram_w16_l1024_id0_1_1_wdata;
        ram_w16_l1024_id0_1_1_rdata_out <= ram_w16_l1024_id0_1_1_wdata;
      end else begin
        ram_w16_l1024_id0_1_1_rdata_out <= mem[ram_w16_l1024_id0_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id1_0
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id1_0_0_addr,
  output [16-1:0] ram_w16_l1024_id1_0_0_rdata,
  input [16-1:0] ram_w16_l1024_id1_0_0_wdata,
  input ram_w16_l1024_id1_0_0_wenable,
  input ram_w16_l1024_id1_0_0_enable,
  input [9-1:0] ram_w16_l1024_id1_0_1_addr,
  output [16-1:0] ram_w16_l1024_id1_0_1_rdata,
  input [16-1:0] ram_w16_l1024_id1_0_1_wdata,
  input ram_w16_l1024_id1_0_1_wenable,
  input ram_w16_l1024_id1_0_1_enable
);

  reg [16-1:0] ram_w16_l1024_id1_0_0_rdata_out;
  assign ram_w16_l1024_id1_0_0_rdata = ram_w16_l1024_id1_0_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id1_0_1_rdata_out;
  assign ram_w16_l1024_id1_0_1_rdata = ram_w16_l1024_id1_0_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id1_0_0_enable) begin
      if(ram_w16_l1024_id1_0_0_wenable) begin
        mem[ram_w16_l1024_id1_0_0_addr] <= ram_w16_l1024_id1_0_0_wdata;
        ram_w16_l1024_id1_0_0_rdata_out <= ram_w16_l1024_id1_0_0_wdata;
      end else begin
        ram_w16_l1024_id1_0_0_rdata_out <= mem[ram_w16_l1024_id1_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id1_0_1_enable) begin
      if(ram_w16_l1024_id1_0_1_wenable) begin
        mem[ram_w16_l1024_id1_0_1_addr] <= ram_w16_l1024_id1_0_1_wdata;
        ram_w16_l1024_id1_0_1_rdata_out <= ram_w16_l1024_id1_0_1_wdata;
      end else begin
        ram_w16_l1024_id1_0_1_rdata_out <= mem[ram_w16_l1024_id1_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id1_1
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id1_1_0_addr,
  output [16-1:0] ram_w16_l1024_id1_1_0_rdata,
  input [16-1:0] ram_w16_l1024_id1_1_0_wdata,
  input ram_w16_l1024_id1_1_0_wenable,
  input ram_w16_l1024_id1_1_0_enable,
  input [9-1:0] ram_w16_l1024_id1_1_1_addr,
  output [16-1:0] ram_w16_l1024_id1_1_1_rdata,
  input [16-1:0] ram_w16_l1024_id1_1_1_wdata,
  input ram_w16_l1024_id1_1_1_wenable,
  input ram_w16_l1024_id1_1_1_enable
);

  reg [16-1:0] ram_w16_l1024_id1_1_0_rdata_out;
  assign ram_w16_l1024_id1_1_0_rdata = ram_w16_l1024_id1_1_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id1_1_1_rdata_out;
  assign ram_w16_l1024_id1_1_1_rdata = ram_w16_l1024_id1_1_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id1_1_0_enable) begin
      if(ram_w16_l1024_id1_1_0_wenable) begin
        mem[ram_w16_l1024_id1_1_0_addr] <= ram_w16_l1024_id1_1_0_wdata;
        ram_w16_l1024_id1_1_0_rdata_out <= ram_w16_l1024_id1_1_0_wdata;
      end else begin
        ram_w16_l1024_id1_1_0_rdata_out <= mem[ram_w16_l1024_id1_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id1_1_1_enable) begin
      if(ram_w16_l1024_id1_1_1_wenable) begin
        mem[ram_w16_l1024_id1_1_1_addr] <= ram_w16_l1024_id1_1_1_wdata;
        ram_w16_l1024_id1_1_1_rdata_out <= ram_w16_l1024_id1_1_1_wdata;
      end else begin
        ram_w16_l1024_id1_1_1_rdata_out <= mem[ram_w16_l1024_id1_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id2_0
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id2_0_0_addr,
  output [16-1:0] ram_w16_l1024_id2_0_0_rdata,
  input [16-1:0] ram_w16_l1024_id2_0_0_wdata,
  input ram_w16_l1024_id2_0_0_wenable,
  input ram_w16_l1024_id2_0_0_enable,
  input [9-1:0] ram_w16_l1024_id2_0_1_addr,
  output [16-1:0] ram_w16_l1024_id2_0_1_rdata,
  input [16-1:0] ram_w16_l1024_id2_0_1_wdata,
  input ram_w16_l1024_id2_0_1_wenable,
  input ram_w16_l1024_id2_0_1_enable
);

  reg [16-1:0] ram_w16_l1024_id2_0_0_rdata_out;
  assign ram_w16_l1024_id2_0_0_rdata = ram_w16_l1024_id2_0_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id2_0_1_rdata_out;
  assign ram_w16_l1024_id2_0_1_rdata = ram_w16_l1024_id2_0_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id2_0_0_enable) begin
      if(ram_w16_l1024_id2_0_0_wenable) begin
        mem[ram_w16_l1024_id2_0_0_addr] <= ram_w16_l1024_id2_0_0_wdata;
        ram_w16_l1024_id2_0_0_rdata_out <= ram_w16_l1024_id2_0_0_wdata;
      end else begin
        ram_w16_l1024_id2_0_0_rdata_out <= mem[ram_w16_l1024_id2_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id2_0_1_enable) begin
      if(ram_w16_l1024_id2_0_1_wenable) begin
        mem[ram_w16_l1024_id2_0_1_addr] <= ram_w16_l1024_id2_0_1_wdata;
        ram_w16_l1024_id2_0_1_rdata_out <= ram_w16_l1024_id2_0_1_wdata;
      end else begin
        ram_w16_l1024_id2_0_1_rdata_out <= mem[ram_w16_l1024_id2_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id2_1
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id2_1_0_addr,
  output [16-1:0] ram_w16_l1024_id2_1_0_rdata,
  input [16-1:0] ram_w16_l1024_id2_1_0_wdata,
  input ram_w16_l1024_id2_1_0_wenable,
  input ram_w16_l1024_id2_1_0_enable,
  input [9-1:0] ram_w16_l1024_id2_1_1_addr,
  output [16-1:0] ram_w16_l1024_id2_1_1_rdata,
  input [16-1:0] ram_w16_l1024_id2_1_1_wdata,
  input ram_w16_l1024_id2_1_1_wenable,
  input ram_w16_l1024_id2_1_1_enable
);

  reg [16-1:0] ram_w16_l1024_id2_1_0_rdata_out;
  assign ram_w16_l1024_id2_1_0_rdata = ram_w16_l1024_id2_1_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id2_1_1_rdata_out;
  assign ram_w16_l1024_id2_1_1_rdata = ram_w16_l1024_id2_1_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id2_1_0_enable) begin
      if(ram_w16_l1024_id2_1_0_wenable) begin
        mem[ram_w16_l1024_id2_1_0_addr] <= ram_w16_l1024_id2_1_0_wdata;
        ram_w16_l1024_id2_1_0_rdata_out <= ram_w16_l1024_id2_1_0_wdata;
      end else begin
        ram_w16_l1024_id2_1_0_rdata_out <= mem[ram_w16_l1024_id2_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id2_1_1_enable) begin
      if(ram_w16_l1024_id2_1_1_wenable) begin
        mem[ram_w16_l1024_id2_1_1_addr] <= ram_w16_l1024_id2_1_1_wdata;
        ram_w16_l1024_id2_1_1_rdata_out <= ram_w16_l1024_id2_1_1_wdata;
      end else begin
        ram_w16_l1024_id2_1_1_rdata_out <= mem[ram_w16_l1024_id2_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id3_0
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id3_0_0_addr,
  output [16-1:0] ram_w16_l1024_id3_0_0_rdata,
  input [16-1:0] ram_w16_l1024_id3_0_0_wdata,
  input ram_w16_l1024_id3_0_0_wenable,
  input ram_w16_l1024_id3_0_0_enable,
  input [9-1:0] ram_w16_l1024_id3_0_1_addr,
  output [16-1:0] ram_w16_l1024_id3_0_1_rdata,
  input [16-1:0] ram_w16_l1024_id3_0_1_wdata,
  input ram_w16_l1024_id3_0_1_wenable,
  input ram_w16_l1024_id3_0_1_enable
);

  reg [16-1:0] ram_w16_l1024_id3_0_0_rdata_out;
  assign ram_w16_l1024_id3_0_0_rdata = ram_w16_l1024_id3_0_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id3_0_1_rdata_out;
  assign ram_w16_l1024_id3_0_1_rdata = ram_w16_l1024_id3_0_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id3_0_0_enable) begin
      if(ram_w16_l1024_id3_0_0_wenable) begin
        mem[ram_w16_l1024_id3_0_0_addr] <= ram_w16_l1024_id3_0_0_wdata;
        ram_w16_l1024_id3_0_0_rdata_out <= ram_w16_l1024_id3_0_0_wdata;
      end else begin
        ram_w16_l1024_id3_0_0_rdata_out <= mem[ram_w16_l1024_id3_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id3_0_1_enable) begin
      if(ram_w16_l1024_id3_0_1_wenable) begin
        mem[ram_w16_l1024_id3_0_1_addr] <= ram_w16_l1024_id3_0_1_wdata;
        ram_w16_l1024_id3_0_1_rdata_out <= ram_w16_l1024_id3_0_1_wdata;
      end else begin
        ram_w16_l1024_id3_0_1_rdata_out <= mem[ram_w16_l1024_id3_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id3_1
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id3_1_0_addr,
  output [16-1:0] ram_w16_l1024_id3_1_0_rdata,
  input [16-1:0] ram_w16_l1024_id3_1_0_wdata,
  input ram_w16_l1024_id3_1_0_wenable,
  input ram_w16_l1024_id3_1_0_enable,
  input [9-1:0] ram_w16_l1024_id3_1_1_addr,
  output [16-1:0] ram_w16_l1024_id3_1_1_rdata,
  input [16-1:0] ram_w16_l1024_id3_1_1_wdata,
  input ram_w16_l1024_id3_1_1_wenable,
  input ram_w16_l1024_id3_1_1_enable
);

  reg [16-1:0] ram_w16_l1024_id3_1_0_rdata_out;
  assign ram_w16_l1024_id3_1_0_rdata = ram_w16_l1024_id3_1_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id3_1_1_rdata_out;
  assign ram_w16_l1024_id3_1_1_rdata = ram_w16_l1024_id3_1_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id3_1_0_enable) begin
      if(ram_w16_l1024_id3_1_0_wenable) begin
        mem[ram_w16_l1024_id3_1_0_addr] <= ram_w16_l1024_id3_1_0_wdata;
        ram_w16_l1024_id3_1_0_rdata_out <= ram_w16_l1024_id3_1_0_wdata;
      end else begin
        ram_w16_l1024_id3_1_0_rdata_out <= mem[ram_w16_l1024_id3_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id3_1_1_enable) begin
      if(ram_w16_l1024_id3_1_1_wenable) begin
        mem[ram_w16_l1024_id3_1_1_addr] <= ram_w16_l1024_id3_1_1_wdata;
        ram_w16_l1024_id3_1_1_rdata_out <= ram_w16_l1024_id3_1_1_wdata;
      end else begin
        ram_w16_l1024_id3_1_1_rdata_out <= mem[ram_w16_l1024_id3_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id4_0
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id4_0_0_addr,
  output [16-1:0] ram_w16_l1024_id4_0_0_rdata,
  input [16-1:0] ram_w16_l1024_id4_0_0_wdata,
  input ram_w16_l1024_id4_0_0_wenable,
  input ram_w16_l1024_id4_0_0_enable,
  input [9-1:0] ram_w16_l1024_id4_0_1_addr,
  output [16-1:0] ram_w16_l1024_id4_0_1_rdata,
  input [16-1:0] ram_w16_l1024_id4_0_1_wdata,
  input ram_w16_l1024_id4_0_1_wenable,
  input ram_w16_l1024_id4_0_1_enable
);

  reg [16-1:0] ram_w16_l1024_id4_0_0_rdata_out;
  assign ram_w16_l1024_id4_0_0_rdata = ram_w16_l1024_id4_0_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id4_0_1_rdata_out;
  assign ram_w16_l1024_id4_0_1_rdata = ram_w16_l1024_id4_0_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id4_0_0_enable) begin
      if(ram_w16_l1024_id4_0_0_wenable) begin
        mem[ram_w16_l1024_id4_0_0_addr] <= ram_w16_l1024_id4_0_0_wdata;
        ram_w16_l1024_id4_0_0_rdata_out <= ram_w16_l1024_id4_0_0_wdata;
      end else begin
        ram_w16_l1024_id4_0_0_rdata_out <= mem[ram_w16_l1024_id4_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id4_0_1_enable) begin
      if(ram_w16_l1024_id4_0_1_wenable) begin
        mem[ram_w16_l1024_id4_0_1_addr] <= ram_w16_l1024_id4_0_1_wdata;
        ram_w16_l1024_id4_0_1_rdata_out <= ram_w16_l1024_id4_0_1_wdata;
      end else begin
        ram_w16_l1024_id4_0_1_rdata_out <= mem[ram_w16_l1024_id4_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id4_1
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id4_1_0_addr,
  output [16-1:0] ram_w16_l1024_id4_1_0_rdata,
  input [16-1:0] ram_w16_l1024_id4_1_0_wdata,
  input ram_w16_l1024_id4_1_0_wenable,
  input ram_w16_l1024_id4_1_0_enable,
  input [9-1:0] ram_w16_l1024_id4_1_1_addr,
  output [16-1:0] ram_w16_l1024_id4_1_1_rdata,
  input [16-1:0] ram_w16_l1024_id4_1_1_wdata,
  input ram_w16_l1024_id4_1_1_wenable,
  input ram_w16_l1024_id4_1_1_enable
);

  reg [16-1:0] ram_w16_l1024_id4_1_0_rdata_out;
  assign ram_w16_l1024_id4_1_0_rdata = ram_w16_l1024_id4_1_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id4_1_1_rdata_out;
  assign ram_w16_l1024_id4_1_1_rdata = ram_w16_l1024_id4_1_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id4_1_0_enable) begin
      if(ram_w16_l1024_id4_1_0_wenable) begin
        mem[ram_w16_l1024_id4_1_0_addr] <= ram_w16_l1024_id4_1_0_wdata;
        ram_w16_l1024_id4_1_0_rdata_out <= ram_w16_l1024_id4_1_0_wdata;
      end else begin
        ram_w16_l1024_id4_1_0_rdata_out <= mem[ram_w16_l1024_id4_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id4_1_1_enable) begin
      if(ram_w16_l1024_id4_1_1_wenable) begin
        mem[ram_w16_l1024_id4_1_1_addr] <= ram_w16_l1024_id4_1_1_wdata;
        ram_w16_l1024_id4_1_1_rdata_out <= ram_w16_l1024_id4_1_1_wdata;
      end else begin
        ram_w16_l1024_id4_1_1_rdata_out <= mem[ram_w16_l1024_id4_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id5_0
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id5_0_0_addr,
  output [16-1:0] ram_w16_l1024_id5_0_0_rdata,
  input [16-1:0] ram_w16_l1024_id5_0_0_wdata,
  input ram_w16_l1024_id5_0_0_wenable,
  input ram_w16_l1024_id5_0_0_enable,
  input [9-1:0] ram_w16_l1024_id5_0_1_addr,
  output [16-1:0] ram_w16_l1024_id5_0_1_rdata,
  input [16-1:0] ram_w16_l1024_id5_0_1_wdata,
  input ram_w16_l1024_id5_0_1_wenable,
  input ram_w16_l1024_id5_0_1_enable
);

  reg [16-1:0] ram_w16_l1024_id5_0_0_rdata_out;
  assign ram_w16_l1024_id5_0_0_rdata = ram_w16_l1024_id5_0_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id5_0_1_rdata_out;
  assign ram_w16_l1024_id5_0_1_rdata = ram_w16_l1024_id5_0_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id5_0_0_enable) begin
      if(ram_w16_l1024_id5_0_0_wenable) begin
        mem[ram_w16_l1024_id5_0_0_addr] <= ram_w16_l1024_id5_0_0_wdata;
        ram_w16_l1024_id5_0_0_rdata_out <= ram_w16_l1024_id5_0_0_wdata;
      end else begin
        ram_w16_l1024_id5_0_0_rdata_out <= mem[ram_w16_l1024_id5_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id5_0_1_enable) begin
      if(ram_w16_l1024_id5_0_1_wenable) begin
        mem[ram_w16_l1024_id5_0_1_addr] <= ram_w16_l1024_id5_0_1_wdata;
        ram_w16_l1024_id5_0_1_rdata_out <= ram_w16_l1024_id5_0_1_wdata;
      end else begin
        ram_w16_l1024_id5_0_1_rdata_out <= mem[ram_w16_l1024_id5_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id5_1
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id5_1_0_addr,
  output [16-1:0] ram_w16_l1024_id5_1_0_rdata,
  input [16-1:0] ram_w16_l1024_id5_1_0_wdata,
  input ram_w16_l1024_id5_1_0_wenable,
  input ram_w16_l1024_id5_1_0_enable,
  input [9-1:0] ram_w16_l1024_id5_1_1_addr,
  output [16-1:0] ram_w16_l1024_id5_1_1_rdata,
  input [16-1:0] ram_w16_l1024_id5_1_1_wdata,
  input ram_w16_l1024_id5_1_1_wenable,
  input ram_w16_l1024_id5_1_1_enable
);

  reg [16-1:0] ram_w16_l1024_id5_1_0_rdata_out;
  assign ram_w16_l1024_id5_1_0_rdata = ram_w16_l1024_id5_1_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id5_1_1_rdata_out;
  assign ram_w16_l1024_id5_1_1_rdata = ram_w16_l1024_id5_1_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id5_1_0_enable) begin
      if(ram_w16_l1024_id5_1_0_wenable) begin
        mem[ram_w16_l1024_id5_1_0_addr] <= ram_w16_l1024_id5_1_0_wdata;
        ram_w16_l1024_id5_1_0_rdata_out <= ram_w16_l1024_id5_1_0_wdata;
      end else begin
        ram_w16_l1024_id5_1_0_rdata_out <= mem[ram_w16_l1024_id5_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id5_1_1_enable) begin
      if(ram_w16_l1024_id5_1_1_wenable) begin
        mem[ram_w16_l1024_id5_1_1_addr] <= ram_w16_l1024_id5_1_1_wdata;
        ram_w16_l1024_id5_1_1_rdata_out <= ram_w16_l1024_id5_1_1_wdata;
      end else begin
        ram_w16_l1024_id5_1_1_rdata_out <= mem[ram_w16_l1024_id5_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id6_0
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id6_0_0_addr,
  output [16-1:0] ram_w16_l1024_id6_0_0_rdata,
  input [16-1:0] ram_w16_l1024_id6_0_0_wdata,
  input ram_w16_l1024_id6_0_0_wenable,
  input ram_w16_l1024_id6_0_0_enable,
  input [9-1:0] ram_w16_l1024_id6_0_1_addr,
  output [16-1:0] ram_w16_l1024_id6_0_1_rdata,
  input [16-1:0] ram_w16_l1024_id6_0_1_wdata,
  input ram_w16_l1024_id6_0_1_wenable,
  input ram_w16_l1024_id6_0_1_enable
);

  reg [16-1:0] ram_w16_l1024_id6_0_0_rdata_out;
  assign ram_w16_l1024_id6_0_0_rdata = ram_w16_l1024_id6_0_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id6_0_1_rdata_out;
  assign ram_w16_l1024_id6_0_1_rdata = ram_w16_l1024_id6_0_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id6_0_0_enable) begin
      if(ram_w16_l1024_id6_0_0_wenable) begin
        mem[ram_w16_l1024_id6_0_0_addr] <= ram_w16_l1024_id6_0_0_wdata;
        ram_w16_l1024_id6_0_0_rdata_out <= ram_w16_l1024_id6_0_0_wdata;
      end else begin
        ram_w16_l1024_id6_0_0_rdata_out <= mem[ram_w16_l1024_id6_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id6_0_1_enable) begin
      if(ram_w16_l1024_id6_0_1_wenable) begin
        mem[ram_w16_l1024_id6_0_1_addr] <= ram_w16_l1024_id6_0_1_wdata;
        ram_w16_l1024_id6_0_1_rdata_out <= ram_w16_l1024_id6_0_1_wdata;
      end else begin
        ram_w16_l1024_id6_0_1_rdata_out <= mem[ram_w16_l1024_id6_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id6_1
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id6_1_0_addr,
  output [16-1:0] ram_w16_l1024_id6_1_0_rdata,
  input [16-1:0] ram_w16_l1024_id6_1_0_wdata,
  input ram_w16_l1024_id6_1_0_wenable,
  input ram_w16_l1024_id6_1_0_enable,
  input [9-1:0] ram_w16_l1024_id6_1_1_addr,
  output [16-1:0] ram_w16_l1024_id6_1_1_rdata,
  input [16-1:0] ram_w16_l1024_id6_1_1_wdata,
  input ram_w16_l1024_id6_1_1_wenable,
  input ram_w16_l1024_id6_1_1_enable
);

  reg [16-1:0] ram_w16_l1024_id6_1_0_rdata_out;
  assign ram_w16_l1024_id6_1_0_rdata = ram_w16_l1024_id6_1_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id6_1_1_rdata_out;
  assign ram_w16_l1024_id6_1_1_rdata = ram_w16_l1024_id6_1_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id6_1_0_enable) begin
      if(ram_w16_l1024_id6_1_0_wenable) begin
        mem[ram_w16_l1024_id6_1_0_addr] <= ram_w16_l1024_id6_1_0_wdata;
        ram_w16_l1024_id6_1_0_rdata_out <= ram_w16_l1024_id6_1_0_wdata;
      end else begin
        ram_w16_l1024_id6_1_0_rdata_out <= mem[ram_w16_l1024_id6_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id6_1_1_enable) begin
      if(ram_w16_l1024_id6_1_1_wenable) begin
        mem[ram_w16_l1024_id6_1_1_addr] <= ram_w16_l1024_id6_1_1_wdata;
        ram_w16_l1024_id6_1_1_rdata_out <= ram_w16_l1024_id6_1_1_wdata;
      end else begin
        ram_w16_l1024_id6_1_1_rdata_out <= mem[ram_w16_l1024_id6_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id7_0
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id7_0_0_addr,
  output [16-1:0] ram_w16_l1024_id7_0_0_rdata,
  input [16-1:0] ram_w16_l1024_id7_0_0_wdata,
  input ram_w16_l1024_id7_0_0_wenable,
  input ram_w16_l1024_id7_0_0_enable,
  input [9-1:0] ram_w16_l1024_id7_0_1_addr,
  output [16-1:0] ram_w16_l1024_id7_0_1_rdata,
  input [16-1:0] ram_w16_l1024_id7_0_1_wdata,
  input ram_w16_l1024_id7_0_1_wenable,
  input ram_w16_l1024_id7_0_1_enable
);

  reg [16-1:0] ram_w16_l1024_id7_0_0_rdata_out;
  assign ram_w16_l1024_id7_0_0_rdata = ram_w16_l1024_id7_0_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id7_0_1_rdata_out;
  assign ram_w16_l1024_id7_0_1_rdata = ram_w16_l1024_id7_0_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id7_0_0_enable) begin
      if(ram_w16_l1024_id7_0_0_wenable) begin
        mem[ram_w16_l1024_id7_0_0_addr] <= ram_w16_l1024_id7_0_0_wdata;
        ram_w16_l1024_id7_0_0_rdata_out <= ram_w16_l1024_id7_0_0_wdata;
      end else begin
        ram_w16_l1024_id7_0_0_rdata_out <= mem[ram_w16_l1024_id7_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id7_0_1_enable) begin
      if(ram_w16_l1024_id7_0_1_wenable) begin
        mem[ram_w16_l1024_id7_0_1_addr] <= ram_w16_l1024_id7_0_1_wdata;
        ram_w16_l1024_id7_0_1_rdata_out <= ram_w16_l1024_id7_0_1_wdata;
      end else begin
        ram_w16_l1024_id7_0_1_rdata_out <= mem[ram_w16_l1024_id7_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id7_1
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id7_1_0_addr,
  output [16-1:0] ram_w16_l1024_id7_1_0_rdata,
  input [16-1:0] ram_w16_l1024_id7_1_0_wdata,
  input ram_w16_l1024_id7_1_0_wenable,
  input ram_w16_l1024_id7_1_0_enable,
  input [9-1:0] ram_w16_l1024_id7_1_1_addr,
  output [16-1:0] ram_w16_l1024_id7_1_1_rdata,
  input [16-1:0] ram_w16_l1024_id7_1_1_wdata,
  input ram_w16_l1024_id7_1_1_wenable,
  input ram_w16_l1024_id7_1_1_enable
);

  reg [16-1:0] ram_w16_l1024_id7_1_0_rdata_out;
  assign ram_w16_l1024_id7_1_0_rdata = ram_w16_l1024_id7_1_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id7_1_1_rdata_out;
  assign ram_w16_l1024_id7_1_1_rdata = ram_w16_l1024_id7_1_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id7_1_0_enable) begin
      if(ram_w16_l1024_id7_1_0_wenable) begin
        mem[ram_w16_l1024_id7_1_0_addr] <= ram_w16_l1024_id7_1_0_wdata;
        ram_w16_l1024_id7_1_0_rdata_out <= ram_w16_l1024_id7_1_0_wdata;
      end else begin
        ram_w16_l1024_id7_1_0_rdata_out <= mem[ram_w16_l1024_id7_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id7_1_1_enable) begin
      if(ram_w16_l1024_id7_1_1_wenable) begin
        mem[ram_w16_l1024_id7_1_1_addr] <= ram_w16_l1024_id7_1_1_wdata;
        ram_w16_l1024_id7_1_1_rdata_out <= ram_w16_l1024_id7_1_1_wdata;
      end else begin
        ram_w16_l1024_id7_1_1_rdata_out <= mem[ram_w16_l1024_id7_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id8_0
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id8_0_0_addr,
  output [16-1:0] ram_w16_l1024_id8_0_0_rdata,
  input [16-1:0] ram_w16_l1024_id8_0_0_wdata,
  input ram_w16_l1024_id8_0_0_wenable,
  input ram_w16_l1024_id8_0_0_enable,
  input [9-1:0] ram_w16_l1024_id8_0_1_addr,
  output [16-1:0] ram_w16_l1024_id8_0_1_rdata,
  input [16-1:0] ram_w16_l1024_id8_0_1_wdata,
  input ram_w16_l1024_id8_0_1_wenable,
  input ram_w16_l1024_id8_0_1_enable
);

  reg [16-1:0] ram_w16_l1024_id8_0_0_rdata_out;
  assign ram_w16_l1024_id8_0_0_rdata = ram_w16_l1024_id8_0_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id8_0_1_rdata_out;
  assign ram_w16_l1024_id8_0_1_rdata = ram_w16_l1024_id8_0_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id8_0_0_enable) begin
      if(ram_w16_l1024_id8_0_0_wenable) begin
        mem[ram_w16_l1024_id8_0_0_addr] <= ram_w16_l1024_id8_0_0_wdata;
        ram_w16_l1024_id8_0_0_rdata_out <= ram_w16_l1024_id8_0_0_wdata;
      end else begin
        ram_w16_l1024_id8_0_0_rdata_out <= mem[ram_w16_l1024_id8_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id8_0_1_enable) begin
      if(ram_w16_l1024_id8_0_1_wenable) begin
        mem[ram_w16_l1024_id8_0_1_addr] <= ram_w16_l1024_id8_0_1_wdata;
        ram_w16_l1024_id8_0_1_rdata_out <= ram_w16_l1024_id8_0_1_wdata;
      end else begin
        ram_w16_l1024_id8_0_1_rdata_out <= mem[ram_w16_l1024_id8_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id8_1
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id8_1_0_addr,
  output [16-1:0] ram_w16_l1024_id8_1_0_rdata,
  input [16-1:0] ram_w16_l1024_id8_1_0_wdata,
  input ram_w16_l1024_id8_1_0_wenable,
  input ram_w16_l1024_id8_1_0_enable,
  input [9-1:0] ram_w16_l1024_id8_1_1_addr,
  output [16-1:0] ram_w16_l1024_id8_1_1_rdata,
  input [16-1:0] ram_w16_l1024_id8_1_1_wdata,
  input ram_w16_l1024_id8_1_1_wenable,
  input ram_w16_l1024_id8_1_1_enable
);

  reg [16-1:0] ram_w16_l1024_id8_1_0_rdata_out;
  assign ram_w16_l1024_id8_1_0_rdata = ram_w16_l1024_id8_1_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id8_1_1_rdata_out;
  assign ram_w16_l1024_id8_1_1_rdata = ram_w16_l1024_id8_1_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id8_1_0_enable) begin
      if(ram_w16_l1024_id8_1_0_wenable) begin
        mem[ram_w16_l1024_id8_1_0_addr] <= ram_w16_l1024_id8_1_0_wdata;
        ram_w16_l1024_id8_1_0_rdata_out <= ram_w16_l1024_id8_1_0_wdata;
      end else begin
        ram_w16_l1024_id8_1_0_rdata_out <= mem[ram_w16_l1024_id8_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id8_1_1_enable) begin
      if(ram_w16_l1024_id8_1_1_wenable) begin
        mem[ram_w16_l1024_id8_1_1_addr] <= ram_w16_l1024_id8_1_1_wdata;
        ram_w16_l1024_id8_1_1_rdata_out <= ram_w16_l1024_id8_1_1_wdata;
      end else begin
        ram_w16_l1024_id8_1_1_rdata_out <= mem[ram_w16_l1024_id8_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id9_0
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id9_0_0_addr,
  output [16-1:0] ram_w16_l1024_id9_0_0_rdata,
  input [16-1:0] ram_w16_l1024_id9_0_0_wdata,
  input ram_w16_l1024_id9_0_0_wenable,
  input ram_w16_l1024_id9_0_0_enable,
  input [9-1:0] ram_w16_l1024_id9_0_1_addr,
  output [16-1:0] ram_w16_l1024_id9_0_1_rdata,
  input [16-1:0] ram_w16_l1024_id9_0_1_wdata,
  input ram_w16_l1024_id9_0_1_wenable,
  input ram_w16_l1024_id9_0_1_enable
);

  reg [16-1:0] ram_w16_l1024_id9_0_0_rdata_out;
  assign ram_w16_l1024_id9_0_0_rdata = ram_w16_l1024_id9_0_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id9_0_1_rdata_out;
  assign ram_w16_l1024_id9_0_1_rdata = ram_w16_l1024_id9_0_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id9_0_0_enable) begin
      if(ram_w16_l1024_id9_0_0_wenable) begin
        mem[ram_w16_l1024_id9_0_0_addr] <= ram_w16_l1024_id9_0_0_wdata;
        ram_w16_l1024_id9_0_0_rdata_out <= ram_w16_l1024_id9_0_0_wdata;
      end else begin
        ram_w16_l1024_id9_0_0_rdata_out <= mem[ram_w16_l1024_id9_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id9_0_1_enable) begin
      if(ram_w16_l1024_id9_0_1_wenable) begin
        mem[ram_w16_l1024_id9_0_1_addr] <= ram_w16_l1024_id9_0_1_wdata;
        ram_w16_l1024_id9_0_1_rdata_out <= ram_w16_l1024_id9_0_1_wdata;
      end else begin
        ram_w16_l1024_id9_0_1_rdata_out <= mem[ram_w16_l1024_id9_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id9_1
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id9_1_0_addr,
  output [16-1:0] ram_w16_l1024_id9_1_0_rdata,
  input [16-1:0] ram_w16_l1024_id9_1_0_wdata,
  input ram_w16_l1024_id9_1_0_wenable,
  input ram_w16_l1024_id9_1_0_enable,
  input [9-1:0] ram_w16_l1024_id9_1_1_addr,
  output [16-1:0] ram_w16_l1024_id9_1_1_rdata,
  input [16-1:0] ram_w16_l1024_id9_1_1_wdata,
  input ram_w16_l1024_id9_1_1_wenable,
  input ram_w16_l1024_id9_1_1_enable
);

  reg [16-1:0] ram_w16_l1024_id9_1_0_rdata_out;
  assign ram_w16_l1024_id9_1_0_rdata = ram_w16_l1024_id9_1_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id9_1_1_rdata_out;
  assign ram_w16_l1024_id9_1_1_rdata = ram_w16_l1024_id9_1_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id9_1_0_enable) begin
      if(ram_w16_l1024_id9_1_0_wenable) begin
        mem[ram_w16_l1024_id9_1_0_addr] <= ram_w16_l1024_id9_1_0_wdata;
        ram_w16_l1024_id9_1_0_rdata_out <= ram_w16_l1024_id9_1_0_wdata;
      end else begin
        ram_w16_l1024_id9_1_0_rdata_out <= mem[ram_w16_l1024_id9_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id9_1_1_enable) begin
      if(ram_w16_l1024_id9_1_1_wenable) begin
        mem[ram_w16_l1024_id9_1_1_addr] <= ram_w16_l1024_id9_1_1_wdata;
        ram_w16_l1024_id9_1_1_rdata_out <= ram_w16_l1024_id9_1_1_wdata;
      end else begin
        ram_w16_l1024_id9_1_1_rdata_out <= mem[ram_w16_l1024_id9_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id10_0
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id10_0_0_addr,
  output [16-1:0] ram_w16_l1024_id10_0_0_rdata,
  input [16-1:0] ram_w16_l1024_id10_0_0_wdata,
  input ram_w16_l1024_id10_0_0_wenable,
  input ram_w16_l1024_id10_0_0_enable,
  input [9-1:0] ram_w16_l1024_id10_0_1_addr,
  output [16-1:0] ram_w16_l1024_id10_0_1_rdata,
  input [16-1:0] ram_w16_l1024_id10_0_1_wdata,
  input ram_w16_l1024_id10_0_1_wenable,
  input ram_w16_l1024_id10_0_1_enable
);

  reg [16-1:0] ram_w16_l1024_id10_0_0_rdata_out;
  assign ram_w16_l1024_id10_0_0_rdata = ram_w16_l1024_id10_0_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id10_0_1_rdata_out;
  assign ram_w16_l1024_id10_0_1_rdata = ram_w16_l1024_id10_0_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id10_0_0_enable) begin
      if(ram_w16_l1024_id10_0_0_wenable) begin
        mem[ram_w16_l1024_id10_0_0_addr] <= ram_w16_l1024_id10_0_0_wdata;
        ram_w16_l1024_id10_0_0_rdata_out <= ram_w16_l1024_id10_0_0_wdata;
      end else begin
        ram_w16_l1024_id10_0_0_rdata_out <= mem[ram_w16_l1024_id10_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id10_0_1_enable) begin
      if(ram_w16_l1024_id10_0_1_wenable) begin
        mem[ram_w16_l1024_id10_0_1_addr] <= ram_w16_l1024_id10_0_1_wdata;
        ram_w16_l1024_id10_0_1_rdata_out <= ram_w16_l1024_id10_0_1_wdata;
      end else begin
        ram_w16_l1024_id10_0_1_rdata_out <= mem[ram_w16_l1024_id10_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l1024_id10_1
(
  input CLK,
  input [9-1:0] ram_w16_l1024_id10_1_0_addr,
  output [16-1:0] ram_w16_l1024_id10_1_0_rdata,
  input [16-1:0] ram_w16_l1024_id10_1_0_wdata,
  input ram_w16_l1024_id10_1_0_wenable,
  input ram_w16_l1024_id10_1_0_enable,
  input [9-1:0] ram_w16_l1024_id10_1_1_addr,
  output [16-1:0] ram_w16_l1024_id10_1_1_rdata,
  input [16-1:0] ram_w16_l1024_id10_1_1_wdata,
  input ram_w16_l1024_id10_1_1_wenable,
  input ram_w16_l1024_id10_1_1_enable
);

  reg [16-1:0] ram_w16_l1024_id10_1_0_rdata_out;
  assign ram_w16_l1024_id10_1_0_rdata = ram_w16_l1024_id10_1_0_rdata_out;
  reg [16-1:0] ram_w16_l1024_id10_1_1_rdata_out;
  assign ram_w16_l1024_id10_1_1_rdata = ram_w16_l1024_id10_1_1_rdata_out;
  reg [16-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w16_l1024_id10_1_0_enable) begin
      if(ram_w16_l1024_id10_1_0_wenable) begin
        mem[ram_w16_l1024_id10_1_0_addr] <= ram_w16_l1024_id10_1_0_wdata;
        ram_w16_l1024_id10_1_0_rdata_out <= ram_w16_l1024_id10_1_0_wdata;
      end else begin
        ram_w16_l1024_id10_1_0_rdata_out <= mem[ram_w16_l1024_id10_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l1024_id10_1_1_enable) begin
      if(ram_w16_l1024_id10_1_1_wenable) begin
        mem[ram_w16_l1024_id10_1_1_addr] <= ram_w16_l1024_id10_1_1_wdata;
        ram_w16_l1024_id10_1_1_rdata_out <= ram_w16_l1024_id10_1_1_wdata;
      end else begin
        ram_w16_l1024_id10_1_1_rdata_out <= mem[ram_w16_l1024_id10_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id0_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id0_0_0_addr,
  output [16-1:0] ram_w16_l512_id0_0_0_rdata,
  input [16-1:0] ram_w16_l512_id0_0_0_wdata,
  input ram_w16_l512_id0_0_0_wenable,
  input ram_w16_l512_id0_0_0_enable,
  input [8-1:0] ram_w16_l512_id0_0_1_addr,
  output [16-1:0] ram_w16_l512_id0_0_1_rdata,
  input [16-1:0] ram_w16_l512_id0_0_1_wdata,
  input ram_w16_l512_id0_0_1_wenable,
  input ram_w16_l512_id0_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id0_0_0_rdata_out;
  assign ram_w16_l512_id0_0_0_rdata = ram_w16_l512_id0_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id0_0_1_rdata_out;
  assign ram_w16_l512_id0_0_1_rdata = ram_w16_l512_id0_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id0_0_0_enable) begin
      if(ram_w16_l512_id0_0_0_wenable) begin
        mem[ram_w16_l512_id0_0_0_addr] <= ram_w16_l512_id0_0_0_wdata;
        ram_w16_l512_id0_0_0_rdata_out <= ram_w16_l512_id0_0_0_wdata;
      end else begin
        ram_w16_l512_id0_0_0_rdata_out <= mem[ram_w16_l512_id0_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id0_0_1_enable) begin
      if(ram_w16_l512_id0_0_1_wenable) begin
        mem[ram_w16_l512_id0_0_1_addr] <= ram_w16_l512_id0_0_1_wdata;
        ram_w16_l512_id0_0_1_rdata_out <= ram_w16_l512_id0_0_1_wdata;
      end else begin
        ram_w16_l512_id0_0_1_rdata_out <= mem[ram_w16_l512_id0_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id0_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id0_1_0_addr,
  output [16-1:0] ram_w16_l512_id0_1_0_rdata,
  input [16-1:0] ram_w16_l512_id0_1_0_wdata,
  input ram_w16_l512_id0_1_0_wenable,
  input ram_w16_l512_id0_1_0_enable,
  input [8-1:0] ram_w16_l512_id0_1_1_addr,
  output [16-1:0] ram_w16_l512_id0_1_1_rdata,
  input [16-1:0] ram_w16_l512_id0_1_1_wdata,
  input ram_w16_l512_id0_1_1_wenable,
  input ram_w16_l512_id0_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id0_1_0_rdata_out;
  assign ram_w16_l512_id0_1_0_rdata = ram_w16_l512_id0_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id0_1_1_rdata_out;
  assign ram_w16_l512_id0_1_1_rdata = ram_w16_l512_id0_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id0_1_0_enable) begin
      if(ram_w16_l512_id0_1_0_wenable) begin
        mem[ram_w16_l512_id0_1_0_addr] <= ram_w16_l512_id0_1_0_wdata;
        ram_w16_l512_id0_1_0_rdata_out <= ram_w16_l512_id0_1_0_wdata;
      end else begin
        ram_w16_l512_id0_1_0_rdata_out <= mem[ram_w16_l512_id0_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id0_1_1_enable) begin
      if(ram_w16_l512_id0_1_1_wenable) begin
        mem[ram_w16_l512_id0_1_1_addr] <= ram_w16_l512_id0_1_1_wdata;
        ram_w16_l512_id0_1_1_rdata_out <= ram_w16_l512_id0_1_1_wdata;
      end else begin
        ram_w16_l512_id0_1_1_rdata_out <= mem[ram_w16_l512_id0_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id1_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id1_0_0_addr,
  output [16-1:0] ram_w16_l512_id1_0_0_rdata,
  input [16-1:0] ram_w16_l512_id1_0_0_wdata,
  input ram_w16_l512_id1_0_0_wenable,
  input ram_w16_l512_id1_0_0_enable,
  input [8-1:0] ram_w16_l512_id1_0_1_addr,
  output [16-1:0] ram_w16_l512_id1_0_1_rdata,
  input [16-1:0] ram_w16_l512_id1_0_1_wdata,
  input ram_w16_l512_id1_0_1_wenable,
  input ram_w16_l512_id1_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id1_0_0_rdata_out;
  assign ram_w16_l512_id1_0_0_rdata = ram_w16_l512_id1_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id1_0_1_rdata_out;
  assign ram_w16_l512_id1_0_1_rdata = ram_w16_l512_id1_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id1_0_0_enable) begin
      if(ram_w16_l512_id1_0_0_wenable) begin
        mem[ram_w16_l512_id1_0_0_addr] <= ram_w16_l512_id1_0_0_wdata;
        ram_w16_l512_id1_0_0_rdata_out <= ram_w16_l512_id1_0_0_wdata;
      end else begin
        ram_w16_l512_id1_0_0_rdata_out <= mem[ram_w16_l512_id1_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id1_0_1_enable) begin
      if(ram_w16_l512_id1_0_1_wenable) begin
        mem[ram_w16_l512_id1_0_1_addr] <= ram_w16_l512_id1_0_1_wdata;
        ram_w16_l512_id1_0_1_rdata_out <= ram_w16_l512_id1_0_1_wdata;
      end else begin
        ram_w16_l512_id1_0_1_rdata_out <= mem[ram_w16_l512_id1_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id1_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id1_1_0_addr,
  output [16-1:0] ram_w16_l512_id1_1_0_rdata,
  input [16-1:0] ram_w16_l512_id1_1_0_wdata,
  input ram_w16_l512_id1_1_0_wenable,
  input ram_w16_l512_id1_1_0_enable,
  input [8-1:0] ram_w16_l512_id1_1_1_addr,
  output [16-1:0] ram_w16_l512_id1_1_1_rdata,
  input [16-1:0] ram_w16_l512_id1_1_1_wdata,
  input ram_w16_l512_id1_1_1_wenable,
  input ram_w16_l512_id1_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id1_1_0_rdata_out;
  assign ram_w16_l512_id1_1_0_rdata = ram_w16_l512_id1_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id1_1_1_rdata_out;
  assign ram_w16_l512_id1_1_1_rdata = ram_w16_l512_id1_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id1_1_0_enable) begin
      if(ram_w16_l512_id1_1_0_wenable) begin
        mem[ram_w16_l512_id1_1_0_addr] <= ram_w16_l512_id1_1_0_wdata;
        ram_w16_l512_id1_1_0_rdata_out <= ram_w16_l512_id1_1_0_wdata;
      end else begin
        ram_w16_l512_id1_1_0_rdata_out <= mem[ram_w16_l512_id1_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id1_1_1_enable) begin
      if(ram_w16_l512_id1_1_1_wenable) begin
        mem[ram_w16_l512_id1_1_1_addr] <= ram_w16_l512_id1_1_1_wdata;
        ram_w16_l512_id1_1_1_rdata_out <= ram_w16_l512_id1_1_1_wdata;
      end else begin
        ram_w16_l512_id1_1_1_rdata_out <= mem[ram_w16_l512_id1_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id2_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id2_0_0_addr,
  output [16-1:0] ram_w16_l512_id2_0_0_rdata,
  input [16-1:0] ram_w16_l512_id2_0_0_wdata,
  input ram_w16_l512_id2_0_0_wenable,
  input ram_w16_l512_id2_0_0_enable,
  input [8-1:0] ram_w16_l512_id2_0_1_addr,
  output [16-1:0] ram_w16_l512_id2_0_1_rdata,
  input [16-1:0] ram_w16_l512_id2_0_1_wdata,
  input ram_w16_l512_id2_0_1_wenable,
  input ram_w16_l512_id2_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id2_0_0_rdata_out;
  assign ram_w16_l512_id2_0_0_rdata = ram_w16_l512_id2_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id2_0_1_rdata_out;
  assign ram_w16_l512_id2_0_1_rdata = ram_w16_l512_id2_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id2_0_0_enable) begin
      if(ram_w16_l512_id2_0_0_wenable) begin
        mem[ram_w16_l512_id2_0_0_addr] <= ram_w16_l512_id2_0_0_wdata;
        ram_w16_l512_id2_0_0_rdata_out <= ram_w16_l512_id2_0_0_wdata;
      end else begin
        ram_w16_l512_id2_0_0_rdata_out <= mem[ram_w16_l512_id2_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id2_0_1_enable) begin
      if(ram_w16_l512_id2_0_1_wenable) begin
        mem[ram_w16_l512_id2_0_1_addr] <= ram_w16_l512_id2_0_1_wdata;
        ram_w16_l512_id2_0_1_rdata_out <= ram_w16_l512_id2_0_1_wdata;
      end else begin
        ram_w16_l512_id2_0_1_rdata_out <= mem[ram_w16_l512_id2_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id2_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id2_1_0_addr,
  output [16-1:0] ram_w16_l512_id2_1_0_rdata,
  input [16-1:0] ram_w16_l512_id2_1_0_wdata,
  input ram_w16_l512_id2_1_0_wenable,
  input ram_w16_l512_id2_1_0_enable,
  input [8-1:0] ram_w16_l512_id2_1_1_addr,
  output [16-1:0] ram_w16_l512_id2_1_1_rdata,
  input [16-1:0] ram_w16_l512_id2_1_1_wdata,
  input ram_w16_l512_id2_1_1_wenable,
  input ram_w16_l512_id2_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id2_1_0_rdata_out;
  assign ram_w16_l512_id2_1_0_rdata = ram_w16_l512_id2_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id2_1_1_rdata_out;
  assign ram_w16_l512_id2_1_1_rdata = ram_w16_l512_id2_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id2_1_0_enable) begin
      if(ram_w16_l512_id2_1_0_wenable) begin
        mem[ram_w16_l512_id2_1_0_addr] <= ram_w16_l512_id2_1_0_wdata;
        ram_w16_l512_id2_1_0_rdata_out <= ram_w16_l512_id2_1_0_wdata;
      end else begin
        ram_w16_l512_id2_1_0_rdata_out <= mem[ram_w16_l512_id2_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id2_1_1_enable) begin
      if(ram_w16_l512_id2_1_1_wenable) begin
        mem[ram_w16_l512_id2_1_1_addr] <= ram_w16_l512_id2_1_1_wdata;
        ram_w16_l512_id2_1_1_rdata_out <= ram_w16_l512_id2_1_1_wdata;
      end else begin
        ram_w16_l512_id2_1_1_rdata_out <= mem[ram_w16_l512_id2_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id3_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id3_0_0_addr,
  output [16-1:0] ram_w16_l512_id3_0_0_rdata,
  input [16-1:0] ram_w16_l512_id3_0_0_wdata,
  input ram_w16_l512_id3_0_0_wenable,
  input ram_w16_l512_id3_0_0_enable,
  input [8-1:0] ram_w16_l512_id3_0_1_addr,
  output [16-1:0] ram_w16_l512_id3_0_1_rdata,
  input [16-1:0] ram_w16_l512_id3_0_1_wdata,
  input ram_w16_l512_id3_0_1_wenable,
  input ram_w16_l512_id3_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id3_0_0_rdata_out;
  assign ram_w16_l512_id3_0_0_rdata = ram_w16_l512_id3_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id3_0_1_rdata_out;
  assign ram_w16_l512_id3_0_1_rdata = ram_w16_l512_id3_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id3_0_0_enable) begin
      if(ram_w16_l512_id3_0_0_wenable) begin
        mem[ram_w16_l512_id3_0_0_addr] <= ram_w16_l512_id3_0_0_wdata;
        ram_w16_l512_id3_0_0_rdata_out <= ram_w16_l512_id3_0_0_wdata;
      end else begin
        ram_w16_l512_id3_0_0_rdata_out <= mem[ram_w16_l512_id3_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id3_0_1_enable) begin
      if(ram_w16_l512_id3_0_1_wenable) begin
        mem[ram_w16_l512_id3_0_1_addr] <= ram_w16_l512_id3_0_1_wdata;
        ram_w16_l512_id3_0_1_rdata_out <= ram_w16_l512_id3_0_1_wdata;
      end else begin
        ram_w16_l512_id3_0_1_rdata_out <= mem[ram_w16_l512_id3_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id3_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id3_1_0_addr,
  output [16-1:0] ram_w16_l512_id3_1_0_rdata,
  input [16-1:0] ram_w16_l512_id3_1_0_wdata,
  input ram_w16_l512_id3_1_0_wenable,
  input ram_w16_l512_id3_1_0_enable,
  input [8-1:0] ram_w16_l512_id3_1_1_addr,
  output [16-1:0] ram_w16_l512_id3_1_1_rdata,
  input [16-1:0] ram_w16_l512_id3_1_1_wdata,
  input ram_w16_l512_id3_1_1_wenable,
  input ram_w16_l512_id3_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id3_1_0_rdata_out;
  assign ram_w16_l512_id3_1_0_rdata = ram_w16_l512_id3_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id3_1_1_rdata_out;
  assign ram_w16_l512_id3_1_1_rdata = ram_w16_l512_id3_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id3_1_0_enable) begin
      if(ram_w16_l512_id3_1_0_wenable) begin
        mem[ram_w16_l512_id3_1_0_addr] <= ram_w16_l512_id3_1_0_wdata;
        ram_w16_l512_id3_1_0_rdata_out <= ram_w16_l512_id3_1_0_wdata;
      end else begin
        ram_w16_l512_id3_1_0_rdata_out <= mem[ram_w16_l512_id3_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id3_1_1_enable) begin
      if(ram_w16_l512_id3_1_1_wenable) begin
        mem[ram_w16_l512_id3_1_1_addr] <= ram_w16_l512_id3_1_1_wdata;
        ram_w16_l512_id3_1_1_rdata_out <= ram_w16_l512_id3_1_1_wdata;
      end else begin
        ram_w16_l512_id3_1_1_rdata_out <= mem[ram_w16_l512_id3_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id4_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id4_0_0_addr,
  output [16-1:0] ram_w16_l512_id4_0_0_rdata,
  input [16-1:0] ram_w16_l512_id4_0_0_wdata,
  input ram_w16_l512_id4_0_0_wenable,
  input ram_w16_l512_id4_0_0_enable,
  input [8-1:0] ram_w16_l512_id4_0_1_addr,
  output [16-1:0] ram_w16_l512_id4_0_1_rdata,
  input [16-1:0] ram_w16_l512_id4_0_1_wdata,
  input ram_w16_l512_id4_0_1_wenable,
  input ram_w16_l512_id4_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id4_0_0_rdata_out;
  assign ram_w16_l512_id4_0_0_rdata = ram_w16_l512_id4_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id4_0_1_rdata_out;
  assign ram_w16_l512_id4_0_1_rdata = ram_w16_l512_id4_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id4_0_0_enable) begin
      if(ram_w16_l512_id4_0_0_wenable) begin
        mem[ram_w16_l512_id4_0_0_addr] <= ram_w16_l512_id4_0_0_wdata;
        ram_w16_l512_id4_0_0_rdata_out <= ram_w16_l512_id4_0_0_wdata;
      end else begin
        ram_w16_l512_id4_0_0_rdata_out <= mem[ram_w16_l512_id4_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id4_0_1_enable) begin
      if(ram_w16_l512_id4_0_1_wenable) begin
        mem[ram_w16_l512_id4_0_1_addr] <= ram_w16_l512_id4_0_1_wdata;
        ram_w16_l512_id4_0_1_rdata_out <= ram_w16_l512_id4_0_1_wdata;
      end else begin
        ram_w16_l512_id4_0_1_rdata_out <= mem[ram_w16_l512_id4_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id4_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id4_1_0_addr,
  output [16-1:0] ram_w16_l512_id4_1_0_rdata,
  input [16-1:0] ram_w16_l512_id4_1_0_wdata,
  input ram_w16_l512_id4_1_0_wenable,
  input ram_w16_l512_id4_1_0_enable,
  input [8-1:0] ram_w16_l512_id4_1_1_addr,
  output [16-1:0] ram_w16_l512_id4_1_1_rdata,
  input [16-1:0] ram_w16_l512_id4_1_1_wdata,
  input ram_w16_l512_id4_1_1_wenable,
  input ram_w16_l512_id4_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id4_1_0_rdata_out;
  assign ram_w16_l512_id4_1_0_rdata = ram_w16_l512_id4_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id4_1_1_rdata_out;
  assign ram_w16_l512_id4_1_1_rdata = ram_w16_l512_id4_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id4_1_0_enable) begin
      if(ram_w16_l512_id4_1_0_wenable) begin
        mem[ram_w16_l512_id4_1_0_addr] <= ram_w16_l512_id4_1_0_wdata;
        ram_w16_l512_id4_1_0_rdata_out <= ram_w16_l512_id4_1_0_wdata;
      end else begin
        ram_w16_l512_id4_1_0_rdata_out <= mem[ram_w16_l512_id4_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id4_1_1_enable) begin
      if(ram_w16_l512_id4_1_1_wenable) begin
        mem[ram_w16_l512_id4_1_1_addr] <= ram_w16_l512_id4_1_1_wdata;
        ram_w16_l512_id4_1_1_rdata_out <= ram_w16_l512_id4_1_1_wdata;
      end else begin
        ram_w16_l512_id4_1_1_rdata_out <= mem[ram_w16_l512_id4_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id5_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id5_0_0_addr,
  output [16-1:0] ram_w16_l512_id5_0_0_rdata,
  input [16-1:0] ram_w16_l512_id5_0_0_wdata,
  input ram_w16_l512_id5_0_0_wenable,
  input ram_w16_l512_id5_0_0_enable,
  input [8-1:0] ram_w16_l512_id5_0_1_addr,
  output [16-1:0] ram_w16_l512_id5_0_1_rdata,
  input [16-1:0] ram_w16_l512_id5_0_1_wdata,
  input ram_w16_l512_id5_0_1_wenable,
  input ram_w16_l512_id5_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id5_0_0_rdata_out;
  assign ram_w16_l512_id5_0_0_rdata = ram_w16_l512_id5_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id5_0_1_rdata_out;
  assign ram_w16_l512_id5_0_1_rdata = ram_w16_l512_id5_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id5_0_0_enable) begin
      if(ram_w16_l512_id5_0_0_wenable) begin
        mem[ram_w16_l512_id5_0_0_addr] <= ram_w16_l512_id5_0_0_wdata;
        ram_w16_l512_id5_0_0_rdata_out <= ram_w16_l512_id5_0_0_wdata;
      end else begin
        ram_w16_l512_id5_0_0_rdata_out <= mem[ram_w16_l512_id5_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id5_0_1_enable) begin
      if(ram_w16_l512_id5_0_1_wenable) begin
        mem[ram_w16_l512_id5_0_1_addr] <= ram_w16_l512_id5_0_1_wdata;
        ram_w16_l512_id5_0_1_rdata_out <= ram_w16_l512_id5_0_1_wdata;
      end else begin
        ram_w16_l512_id5_0_1_rdata_out <= mem[ram_w16_l512_id5_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id5_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id5_1_0_addr,
  output [16-1:0] ram_w16_l512_id5_1_0_rdata,
  input [16-1:0] ram_w16_l512_id5_1_0_wdata,
  input ram_w16_l512_id5_1_0_wenable,
  input ram_w16_l512_id5_1_0_enable,
  input [8-1:0] ram_w16_l512_id5_1_1_addr,
  output [16-1:0] ram_w16_l512_id5_1_1_rdata,
  input [16-1:0] ram_w16_l512_id5_1_1_wdata,
  input ram_w16_l512_id5_1_1_wenable,
  input ram_w16_l512_id5_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id5_1_0_rdata_out;
  assign ram_w16_l512_id5_1_0_rdata = ram_w16_l512_id5_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id5_1_1_rdata_out;
  assign ram_w16_l512_id5_1_1_rdata = ram_w16_l512_id5_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id5_1_0_enable) begin
      if(ram_w16_l512_id5_1_0_wenable) begin
        mem[ram_w16_l512_id5_1_0_addr] <= ram_w16_l512_id5_1_0_wdata;
        ram_w16_l512_id5_1_0_rdata_out <= ram_w16_l512_id5_1_0_wdata;
      end else begin
        ram_w16_l512_id5_1_0_rdata_out <= mem[ram_w16_l512_id5_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id5_1_1_enable) begin
      if(ram_w16_l512_id5_1_1_wenable) begin
        mem[ram_w16_l512_id5_1_1_addr] <= ram_w16_l512_id5_1_1_wdata;
        ram_w16_l512_id5_1_1_rdata_out <= ram_w16_l512_id5_1_1_wdata;
      end else begin
        ram_w16_l512_id5_1_1_rdata_out <= mem[ram_w16_l512_id5_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id6_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id6_0_0_addr,
  output [16-1:0] ram_w16_l512_id6_0_0_rdata,
  input [16-1:0] ram_w16_l512_id6_0_0_wdata,
  input ram_w16_l512_id6_0_0_wenable,
  input ram_w16_l512_id6_0_0_enable,
  input [8-1:0] ram_w16_l512_id6_0_1_addr,
  output [16-1:0] ram_w16_l512_id6_0_1_rdata,
  input [16-1:0] ram_w16_l512_id6_0_1_wdata,
  input ram_w16_l512_id6_0_1_wenable,
  input ram_w16_l512_id6_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id6_0_0_rdata_out;
  assign ram_w16_l512_id6_0_0_rdata = ram_w16_l512_id6_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id6_0_1_rdata_out;
  assign ram_w16_l512_id6_0_1_rdata = ram_w16_l512_id6_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id6_0_0_enable) begin
      if(ram_w16_l512_id6_0_0_wenable) begin
        mem[ram_w16_l512_id6_0_0_addr] <= ram_w16_l512_id6_0_0_wdata;
        ram_w16_l512_id6_0_0_rdata_out <= ram_w16_l512_id6_0_0_wdata;
      end else begin
        ram_w16_l512_id6_0_0_rdata_out <= mem[ram_w16_l512_id6_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id6_0_1_enable) begin
      if(ram_w16_l512_id6_0_1_wenable) begin
        mem[ram_w16_l512_id6_0_1_addr] <= ram_w16_l512_id6_0_1_wdata;
        ram_w16_l512_id6_0_1_rdata_out <= ram_w16_l512_id6_0_1_wdata;
      end else begin
        ram_w16_l512_id6_0_1_rdata_out <= mem[ram_w16_l512_id6_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id6_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id6_1_0_addr,
  output [16-1:0] ram_w16_l512_id6_1_0_rdata,
  input [16-1:0] ram_w16_l512_id6_1_0_wdata,
  input ram_w16_l512_id6_1_0_wenable,
  input ram_w16_l512_id6_1_0_enable,
  input [8-1:0] ram_w16_l512_id6_1_1_addr,
  output [16-1:0] ram_w16_l512_id6_1_1_rdata,
  input [16-1:0] ram_w16_l512_id6_1_1_wdata,
  input ram_w16_l512_id6_1_1_wenable,
  input ram_w16_l512_id6_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id6_1_0_rdata_out;
  assign ram_w16_l512_id6_1_0_rdata = ram_w16_l512_id6_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id6_1_1_rdata_out;
  assign ram_w16_l512_id6_1_1_rdata = ram_w16_l512_id6_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id6_1_0_enable) begin
      if(ram_w16_l512_id6_1_0_wenable) begin
        mem[ram_w16_l512_id6_1_0_addr] <= ram_w16_l512_id6_1_0_wdata;
        ram_w16_l512_id6_1_0_rdata_out <= ram_w16_l512_id6_1_0_wdata;
      end else begin
        ram_w16_l512_id6_1_0_rdata_out <= mem[ram_w16_l512_id6_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id6_1_1_enable) begin
      if(ram_w16_l512_id6_1_1_wenable) begin
        mem[ram_w16_l512_id6_1_1_addr] <= ram_w16_l512_id6_1_1_wdata;
        ram_w16_l512_id6_1_1_rdata_out <= ram_w16_l512_id6_1_1_wdata;
      end else begin
        ram_w16_l512_id6_1_1_rdata_out <= mem[ram_w16_l512_id6_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id7_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id7_0_0_addr,
  output [16-1:0] ram_w16_l512_id7_0_0_rdata,
  input [16-1:0] ram_w16_l512_id7_0_0_wdata,
  input ram_w16_l512_id7_0_0_wenable,
  input ram_w16_l512_id7_0_0_enable,
  input [8-1:0] ram_w16_l512_id7_0_1_addr,
  output [16-1:0] ram_w16_l512_id7_0_1_rdata,
  input [16-1:0] ram_w16_l512_id7_0_1_wdata,
  input ram_w16_l512_id7_0_1_wenable,
  input ram_w16_l512_id7_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id7_0_0_rdata_out;
  assign ram_w16_l512_id7_0_0_rdata = ram_w16_l512_id7_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id7_0_1_rdata_out;
  assign ram_w16_l512_id7_0_1_rdata = ram_w16_l512_id7_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id7_0_0_enable) begin
      if(ram_w16_l512_id7_0_0_wenable) begin
        mem[ram_w16_l512_id7_0_0_addr] <= ram_w16_l512_id7_0_0_wdata;
        ram_w16_l512_id7_0_0_rdata_out <= ram_w16_l512_id7_0_0_wdata;
      end else begin
        ram_w16_l512_id7_0_0_rdata_out <= mem[ram_w16_l512_id7_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id7_0_1_enable) begin
      if(ram_w16_l512_id7_0_1_wenable) begin
        mem[ram_w16_l512_id7_0_1_addr] <= ram_w16_l512_id7_0_1_wdata;
        ram_w16_l512_id7_0_1_rdata_out <= ram_w16_l512_id7_0_1_wdata;
      end else begin
        ram_w16_l512_id7_0_1_rdata_out <= mem[ram_w16_l512_id7_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id7_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id7_1_0_addr,
  output [16-1:0] ram_w16_l512_id7_1_0_rdata,
  input [16-1:0] ram_w16_l512_id7_1_0_wdata,
  input ram_w16_l512_id7_1_0_wenable,
  input ram_w16_l512_id7_1_0_enable,
  input [8-1:0] ram_w16_l512_id7_1_1_addr,
  output [16-1:0] ram_w16_l512_id7_1_1_rdata,
  input [16-1:0] ram_w16_l512_id7_1_1_wdata,
  input ram_w16_l512_id7_1_1_wenable,
  input ram_w16_l512_id7_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id7_1_0_rdata_out;
  assign ram_w16_l512_id7_1_0_rdata = ram_w16_l512_id7_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id7_1_1_rdata_out;
  assign ram_w16_l512_id7_1_1_rdata = ram_w16_l512_id7_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id7_1_0_enable) begin
      if(ram_w16_l512_id7_1_0_wenable) begin
        mem[ram_w16_l512_id7_1_0_addr] <= ram_w16_l512_id7_1_0_wdata;
        ram_w16_l512_id7_1_0_rdata_out <= ram_w16_l512_id7_1_0_wdata;
      end else begin
        ram_w16_l512_id7_1_0_rdata_out <= mem[ram_w16_l512_id7_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id7_1_1_enable) begin
      if(ram_w16_l512_id7_1_1_wenable) begin
        mem[ram_w16_l512_id7_1_1_addr] <= ram_w16_l512_id7_1_1_wdata;
        ram_w16_l512_id7_1_1_rdata_out <= ram_w16_l512_id7_1_1_wdata;
      end else begin
        ram_w16_l512_id7_1_1_rdata_out <= mem[ram_w16_l512_id7_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id8_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id8_0_0_addr,
  output [16-1:0] ram_w16_l512_id8_0_0_rdata,
  input [16-1:0] ram_w16_l512_id8_0_0_wdata,
  input ram_w16_l512_id8_0_0_wenable,
  input ram_w16_l512_id8_0_0_enable,
  input [8-1:0] ram_w16_l512_id8_0_1_addr,
  output [16-1:0] ram_w16_l512_id8_0_1_rdata,
  input [16-1:0] ram_w16_l512_id8_0_1_wdata,
  input ram_w16_l512_id8_0_1_wenable,
  input ram_w16_l512_id8_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id8_0_0_rdata_out;
  assign ram_w16_l512_id8_0_0_rdata = ram_w16_l512_id8_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id8_0_1_rdata_out;
  assign ram_w16_l512_id8_0_1_rdata = ram_w16_l512_id8_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id8_0_0_enable) begin
      if(ram_w16_l512_id8_0_0_wenable) begin
        mem[ram_w16_l512_id8_0_0_addr] <= ram_w16_l512_id8_0_0_wdata;
        ram_w16_l512_id8_0_0_rdata_out <= ram_w16_l512_id8_0_0_wdata;
      end else begin
        ram_w16_l512_id8_0_0_rdata_out <= mem[ram_w16_l512_id8_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id8_0_1_enable) begin
      if(ram_w16_l512_id8_0_1_wenable) begin
        mem[ram_w16_l512_id8_0_1_addr] <= ram_w16_l512_id8_0_1_wdata;
        ram_w16_l512_id8_0_1_rdata_out <= ram_w16_l512_id8_0_1_wdata;
      end else begin
        ram_w16_l512_id8_0_1_rdata_out <= mem[ram_w16_l512_id8_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id8_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id8_1_0_addr,
  output [16-1:0] ram_w16_l512_id8_1_0_rdata,
  input [16-1:0] ram_w16_l512_id8_1_0_wdata,
  input ram_w16_l512_id8_1_0_wenable,
  input ram_w16_l512_id8_1_0_enable,
  input [8-1:0] ram_w16_l512_id8_1_1_addr,
  output [16-1:0] ram_w16_l512_id8_1_1_rdata,
  input [16-1:0] ram_w16_l512_id8_1_1_wdata,
  input ram_w16_l512_id8_1_1_wenable,
  input ram_w16_l512_id8_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id8_1_0_rdata_out;
  assign ram_w16_l512_id8_1_0_rdata = ram_w16_l512_id8_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id8_1_1_rdata_out;
  assign ram_w16_l512_id8_1_1_rdata = ram_w16_l512_id8_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id8_1_0_enable) begin
      if(ram_w16_l512_id8_1_0_wenable) begin
        mem[ram_w16_l512_id8_1_0_addr] <= ram_w16_l512_id8_1_0_wdata;
        ram_w16_l512_id8_1_0_rdata_out <= ram_w16_l512_id8_1_0_wdata;
      end else begin
        ram_w16_l512_id8_1_0_rdata_out <= mem[ram_w16_l512_id8_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id8_1_1_enable) begin
      if(ram_w16_l512_id8_1_1_wenable) begin
        mem[ram_w16_l512_id8_1_1_addr] <= ram_w16_l512_id8_1_1_wdata;
        ram_w16_l512_id8_1_1_rdata_out <= ram_w16_l512_id8_1_1_wdata;
      end else begin
        ram_w16_l512_id8_1_1_rdata_out <= mem[ram_w16_l512_id8_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id9_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id9_0_0_addr,
  output [16-1:0] ram_w16_l512_id9_0_0_rdata,
  input [16-1:0] ram_w16_l512_id9_0_0_wdata,
  input ram_w16_l512_id9_0_0_wenable,
  input ram_w16_l512_id9_0_0_enable,
  input [8-1:0] ram_w16_l512_id9_0_1_addr,
  output [16-1:0] ram_w16_l512_id9_0_1_rdata,
  input [16-1:0] ram_w16_l512_id9_0_1_wdata,
  input ram_w16_l512_id9_0_1_wenable,
  input ram_w16_l512_id9_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id9_0_0_rdata_out;
  assign ram_w16_l512_id9_0_0_rdata = ram_w16_l512_id9_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id9_0_1_rdata_out;
  assign ram_w16_l512_id9_0_1_rdata = ram_w16_l512_id9_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id9_0_0_enable) begin
      if(ram_w16_l512_id9_0_0_wenable) begin
        mem[ram_w16_l512_id9_0_0_addr] <= ram_w16_l512_id9_0_0_wdata;
        ram_w16_l512_id9_0_0_rdata_out <= ram_w16_l512_id9_0_0_wdata;
      end else begin
        ram_w16_l512_id9_0_0_rdata_out <= mem[ram_w16_l512_id9_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id9_0_1_enable) begin
      if(ram_w16_l512_id9_0_1_wenable) begin
        mem[ram_w16_l512_id9_0_1_addr] <= ram_w16_l512_id9_0_1_wdata;
        ram_w16_l512_id9_0_1_rdata_out <= ram_w16_l512_id9_0_1_wdata;
      end else begin
        ram_w16_l512_id9_0_1_rdata_out <= mem[ram_w16_l512_id9_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id9_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id9_1_0_addr,
  output [16-1:0] ram_w16_l512_id9_1_0_rdata,
  input [16-1:0] ram_w16_l512_id9_1_0_wdata,
  input ram_w16_l512_id9_1_0_wenable,
  input ram_w16_l512_id9_1_0_enable,
  input [8-1:0] ram_w16_l512_id9_1_1_addr,
  output [16-1:0] ram_w16_l512_id9_1_1_rdata,
  input [16-1:0] ram_w16_l512_id9_1_1_wdata,
  input ram_w16_l512_id9_1_1_wenable,
  input ram_w16_l512_id9_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id9_1_0_rdata_out;
  assign ram_w16_l512_id9_1_0_rdata = ram_w16_l512_id9_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id9_1_1_rdata_out;
  assign ram_w16_l512_id9_1_1_rdata = ram_w16_l512_id9_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id9_1_0_enable) begin
      if(ram_w16_l512_id9_1_0_wenable) begin
        mem[ram_w16_l512_id9_1_0_addr] <= ram_w16_l512_id9_1_0_wdata;
        ram_w16_l512_id9_1_0_rdata_out <= ram_w16_l512_id9_1_0_wdata;
      end else begin
        ram_w16_l512_id9_1_0_rdata_out <= mem[ram_w16_l512_id9_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id9_1_1_enable) begin
      if(ram_w16_l512_id9_1_1_wenable) begin
        mem[ram_w16_l512_id9_1_1_addr] <= ram_w16_l512_id9_1_1_wdata;
        ram_w16_l512_id9_1_1_rdata_out <= ram_w16_l512_id9_1_1_wdata;
      end else begin
        ram_w16_l512_id9_1_1_rdata_out <= mem[ram_w16_l512_id9_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id10_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id10_0_0_addr,
  output [16-1:0] ram_w16_l512_id10_0_0_rdata,
  input [16-1:0] ram_w16_l512_id10_0_0_wdata,
  input ram_w16_l512_id10_0_0_wenable,
  input ram_w16_l512_id10_0_0_enable,
  input [8-1:0] ram_w16_l512_id10_0_1_addr,
  output [16-1:0] ram_w16_l512_id10_0_1_rdata,
  input [16-1:0] ram_w16_l512_id10_0_1_wdata,
  input ram_w16_l512_id10_0_1_wenable,
  input ram_w16_l512_id10_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id10_0_0_rdata_out;
  assign ram_w16_l512_id10_0_0_rdata = ram_w16_l512_id10_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id10_0_1_rdata_out;
  assign ram_w16_l512_id10_0_1_rdata = ram_w16_l512_id10_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id10_0_0_enable) begin
      if(ram_w16_l512_id10_0_0_wenable) begin
        mem[ram_w16_l512_id10_0_0_addr] <= ram_w16_l512_id10_0_0_wdata;
        ram_w16_l512_id10_0_0_rdata_out <= ram_w16_l512_id10_0_0_wdata;
      end else begin
        ram_w16_l512_id10_0_0_rdata_out <= mem[ram_w16_l512_id10_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id10_0_1_enable) begin
      if(ram_w16_l512_id10_0_1_wenable) begin
        mem[ram_w16_l512_id10_0_1_addr] <= ram_w16_l512_id10_0_1_wdata;
        ram_w16_l512_id10_0_1_rdata_out <= ram_w16_l512_id10_0_1_wdata;
      end else begin
        ram_w16_l512_id10_0_1_rdata_out <= mem[ram_w16_l512_id10_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id10_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id10_1_0_addr,
  output [16-1:0] ram_w16_l512_id10_1_0_rdata,
  input [16-1:0] ram_w16_l512_id10_1_0_wdata,
  input ram_w16_l512_id10_1_0_wenable,
  input ram_w16_l512_id10_1_0_enable,
  input [8-1:0] ram_w16_l512_id10_1_1_addr,
  output [16-1:0] ram_w16_l512_id10_1_1_rdata,
  input [16-1:0] ram_w16_l512_id10_1_1_wdata,
  input ram_w16_l512_id10_1_1_wenable,
  input ram_w16_l512_id10_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id10_1_0_rdata_out;
  assign ram_w16_l512_id10_1_0_rdata = ram_w16_l512_id10_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id10_1_1_rdata_out;
  assign ram_w16_l512_id10_1_1_rdata = ram_w16_l512_id10_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id10_1_0_enable) begin
      if(ram_w16_l512_id10_1_0_wenable) begin
        mem[ram_w16_l512_id10_1_0_addr] <= ram_w16_l512_id10_1_0_wdata;
        ram_w16_l512_id10_1_0_rdata_out <= ram_w16_l512_id10_1_0_wdata;
      end else begin
        ram_w16_l512_id10_1_0_rdata_out <= mem[ram_w16_l512_id10_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id10_1_1_enable) begin
      if(ram_w16_l512_id10_1_1_wenable) begin
        mem[ram_w16_l512_id10_1_1_addr] <= ram_w16_l512_id10_1_1_wdata;
        ram_w16_l512_id10_1_1_rdata_out <= ram_w16_l512_id10_1_1_wdata;
      end else begin
        ram_w16_l512_id10_1_1_rdata_out <= mem[ram_w16_l512_id10_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id11_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id11_0_0_addr,
  output [16-1:0] ram_w16_l512_id11_0_0_rdata,
  input [16-1:0] ram_w16_l512_id11_0_0_wdata,
  input ram_w16_l512_id11_0_0_wenable,
  input ram_w16_l512_id11_0_0_enable,
  input [8-1:0] ram_w16_l512_id11_0_1_addr,
  output [16-1:0] ram_w16_l512_id11_0_1_rdata,
  input [16-1:0] ram_w16_l512_id11_0_1_wdata,
  input ram_w16_l512_id11_0_1_wenable,
  input ram_w16_l512_id11_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id11_0_0_rdata_out;
  assign ram_w16_l512_id11_0_0_rdata = ram_w16_l512_id11_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id11_0_1_rdata_out;
  assign ram_w16_l512_id11_0_1_rdata = ram_w16_l512_id11_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id11_0_0_enable) begin
      if(ram_w16_l512_id11_0_0_wenable) begin
        mem[ram_w16_l512_id11_0_0_addr] <= ram_w16_l512_id11_0_0_wdata;
        ram_w16_l512_id11_0_0_rdata_out <= ram_w16_l512_id11_0_0_wdata;
      end else begin
        ram_w16_l512_id11_0_0_rdata_out <= mem[ram_w16_l512_id11_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id11_0_1_enable) begin
      if(ram_w16_l512_id11_0_1_wenable) begin
        mem[ram_w16_l512_id11_0_1_addr] <= ram_w16_l512_id11_0_1_wdata;
        ram_w16_l512_id11_0_1_rdata_out <= ram_w16_l512_id11_0_1_wdata;
      end else begin
        ram_w16_l512_id11_0_1_rdata_out <= mem[ram_w16_l512_id11_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id11_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id11_1_0_addr,
  output [16-1:0] ram_w16_l512_id11_1_0_rdata,
  input [16-1:0] ram_w16_l512_id11_1_0_wdata,
  input ram_w16_l512_id11_1_0_wenable,
  input ram_w16_l512_id11_1_0_enable,
  input [8-1:0] ram_w16_l512_id11_1_1_addr,
  output [16-1:0] ram_w16_l512_id11_1_1_rdata,
  input [16-1:0] ram_w16_l512_id11_1_1_wdata,
  input ram_w16_l512_id11_1_1_wenable,
  input ram_w16_l512_id11_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id11_1_0_rdata_out;
  assign ram_w16_l512_id11_1_0_rdata = ram_w16_l512_id11_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id11_1_1_rdata_out;
  assign ram_w16_l512_id11_1_1_rdata = ram_w16_l512_id11_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id11_1_0_enable) begin
      if(ram_w16_l512_id11_1_0_wenable) begin
        mem[ram_w16_l512_id11_1_0_addr] <= ram_w16_l512_id11_1_0_wdata;
        ram_w16_l512_id11_1_0_rdata_out <= ram_w16_l512_id11_1_0_wdata;
      end else begin
        ram_w16_l512_id11_1_0_rdata_out <= mem[ram_w16_l512_id11_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id11_1_1_enable) begin
      if(ram_w16_l512_id11_1_1_wenable) begin
        mem[ram_w16_l512_id11_1_1_addr] <= ram_w16_l512_id11_1_1_wdata;
        ram_w16_l512_id11_1_1_rdata_out <= ram_w16_l512_id11_1_1_wdata;
      end else begin
        ram_w16_l512_id11_1_1_rdata_out <= mem[ram_w16_l512_id11_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id12_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id12_0_0_addr,
  output [16-1:0] ram_w16_l512_id12_0_0_rdata,
  input [16-1:0] ram_w16_l512_id12_0_0_wdata,
  input ram_w16_l512_id12_0_0_wenable,
  input ram_w16_l512_id12_0_0_enable,
  input [8-1:0] ram_w16_l512_id12_0_1_addr,
  output [16-1:0] ram_w16_l512_id12_0_1_rdata,
  input [16-1:0] ram_w16_l512_id12_0_1_wdata,
  input ram_w16_l512_id12_0_1_wenable,
  input ram_w16_l512_id12_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id12_0_0_rdata_out;
  assign ram_w16_l512_id12_0_0_rdata = ram_w16_l512_id12_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id12_0_1_rdata_out;
  assign ram_w16_l512_id12_0_1_rdata = ram_w16_l512_id12_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id12_0_0_enable) begin
      if(ram_w16_l512_id12_0_0_wenable) begin
        mem[ram_w16_l512_id12_0_0_addr] <= ram_w16_l512_id12_0_0_wdata;
        ram_w16_l512_id12_0_0_rdata_out <= ram_w16_l512_id12_0_0_wdata;
      end else begin
        ram_w16_l512_id12_0_0_rdata_out <= mem[ram_w16_l512_id12_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id12_0_1_enable) begin
      if(ram_w16_l512_id12_0_1_wenable) begin
        mem[ram_w16_l512_id12_0_1_addr] <= ram_w16_l512_id12_0_1_wdata;
        ram_w16_l512_id12_0_1_rdata_out <= ram_w16_l512_id12_0_1_wdata;
      end else begin
        ram_w16_l512_id12_0_1_rdata_out <= mem[ram_w16_l512_id12_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id12_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id12_1_0_addr,
  output [16-1:0] ram_w16_l512_id12_1_0_rdata,
  input [16-1:0] ram_w16_l512_id12_1_0_wdata,
  input ram_w16_l512_id12_1_0_wenable,
  input ram_w16_l512_id12_1_0_enable,
  input [8-1:0] ram_w16_l512_id12_1_1_addr,
  output [16-1:0] ram_w16_l512_id12_1_1_rdata,
  input [16-1:0] ram_w16_l512_id12_1_1_wdata,
  input ram_w16_l512_id12_1_1_wenable,
  input ram_w16_l512_id12_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id12_1_0_rdata_out;
  assign ram_w16_l512_id12_1_0_rdata = ram_w16_l512_id12_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id12_1_1_rdata_out;
  assign ram_w16_l512_id12_1_1_rdata = ram_w16_l512_id12_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id12_1_0_enable) begin
      if(ram_w16_l512_id12_1_0_wenable) begin
        mem[ram_w16_l512_id12_1_0_addr] <= ram_w16_l512_id12_1_0_wdata;
        ram_w16_l512_id12_1_0_rdata_out <= ram_w16_l512_id12_1_0_wdata;
      end else begin
        ram_w16_l512_id12_1_0_rdata_out <= mem[ram_w16_l512_id12_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id12_1_1_enable) begin
      if(ram_w16_l512_id12_1_1_wenable) begin
        mem[ram_w16_l512_id12_1_1_addr] <= ram_w16_l512_id12_1_1_wdata;
        ram_w16_l512_id12_1_1_rdata_out <= ram_w16_l512_id12_1_1_wdata;
      end else begin
        ram_w16_l512_id12_1_1_rdata_out <= mem[ram_w16_l512_id12_1_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id0
(
  input CLK,
  input [7-1:0] ram_w32_l128_id0_0_addr,
  output [32-1:0] ram_w32_l128_id0_0_rdata,
  input [32-1:0] ram_w32_l128_id0_0_wdata,
  input ram_w32_l128_id0_0_wenable,
  input ram_w32_l128_id0_0_enable,
  input [7-1:0] ram_w32_l128_id0_1_addr,
  output [32-1:0] ram_w32_l128_id0_1_rdata,
  input [32-1:0] ram_w32_l128_id0_1_wdata,
  input ram_w32_l128_id0_1_wenable,
  input ram_w32_l128_id0_1_enable
);

  reg [32-1:0] ram_w32_l128_id0_0_rdata_out;
  assign ram_w32_l128_id0_0_rdata = ram_w32_l128_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id0_1_rdata_out;
  assign ram_w32_l128_id0_1_rdata = ram_w32_l128_id0_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id0_0_enable) begin
      if(ram_w32_l128_id0_0_wenable) begin
        mem[ram_w32_l128_id0_0_addr] <= ram_w32_l128_id0_0_wdata;
        ram_w32_l128_id0_0_rdata_out <= ram_w32_l128_id0_0_wdata;
      end else begin
        ram_w32_l128_id0_0_rdata_out <= mem[ram_w32_l128_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id0_1_enable) begin
      if(ram_w32_l128_id0_1_wenable) begin
        mem[ram_w32_l128_id0_1_addr] <= ram_w32_l128_id0_1_wdata;
        ram_w32_l128_id0_1_rdata_out <= ram_w32_l128_id0_1_wdata;
      end else begin
        ram_w32_l128_id0_1_rdata_out <= mem[ram_w32_l128_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id1
(
  input CLK,
  input [7-1:0] ram_w32_l128_id1_0_addr,
  output [32-1:0] ram_w32_l128_id1_0_rdata,
  input [32-1:0] ram_w32_l128_id1_0_wdata,
  input ram_w32_l128_id1_0_wenable,
  input ram_w32_l128_id1_0_enable,
  input [7-1:0] ram_w32_l128_id1_1_addr,
  output [32-1:0] ram_w32_l128_id1_1_rdata,
  input [32-1:0] ram_w32_l128_id1_1_wdata,
  input ram_w32_l128_id1_1_wenable,
  input ram_w32_l128_id1_1_enable
);

  reg [32-1:0] ram_w32_l128_id1_0_rdata_out;
  assign ram_w32_l128_id1_0_rdata = ram_w32_l128_id1_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id1_1_rdata_out;
  assign ram_w32_l128_id1_1_rdata = ram_w32_l128_id1_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id1_0_enable) begin
      if(ram_w32_l128_id1_0_wenable) begin
        mem[ram_w32_l128_id1_0_addr] <= ram_w32_l128_id1_0_wdata;
        ram_w32_l128_id1_0_rdata_out <= ram_w32_l128_id1_0_wdata;
      end else begin
        ram_w32_l128_id1_0_rdata_out <= mem[ram_w32_l128_id1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id1_1_enable) begin
      if(ram_w32_l128_id1_1_wenable) begin
        mem[ram_w32_l128_id1_1_addr] <= ram_w32_l128_id1_1_wdata;
        ram_w32_l128_id1_1_rdata_out <= ram_w32_l128_id1_1_wdata;
      end else begin
        ram_w32_l128_id1_1_rdata_out <= mem[ram_w32_l128_id1_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id2
(
  input CLK,
  input [7-1:0] ram_w32_l128_id2_0_addr,
  output [32-1:0] ram_w32_l128_id2_0_rdata,
  input [32-1:0] ram_w32_l128_id2_0_wdata,
  input ram_w32_l128_id2_0_wenable,
  input ram_w32_l128_id2_0_enable,
  input [7-1:0] ram_w32_l128_id2_1_addr,
  output [32-1:0] ram_w32_l128_id2_1_rdata,
  input [32-1:0] ram_w32_l128_id2_1_wdata,
  input ram_w32_l128_id2_1_wenable,
  input ram_w32_l128_id2_1_enable
);

  reg [32-1:0] ram_w32_l128_id2_0_rdata_out;
  assign ram_w32_l128_id2_0_rdata = ram_w32_l128_id2_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id2_1_rdata_out;
  assign ram_w32_l128_id2_1_rdata = ram_w32_l128_id2_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id2_0_enable) begin
      if(ram_w32_l128_id2_0_wenable) begin
        mem[ram_w32_l128_id2_0_addr] <= ram_w32_l128_id2_0_wdata;
        ram_w32_l128_id2_0_rdata_out <= ram_w32_l128_id2_0_wdata;
      end else begin
        ram_w32_l128_id2_0_rdata_out <= mem[ram_w32_l128_id2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id2_1_enable) begin
      if(ram_w32_l128_id2_1_wenable) begin
        mem[ram_w32_l128_id2_1_addr] <= ram_w32_l128_id2_1_wdata;
        ram_w32_l128_id2_1_rdata_out <= ram_w32_l128_id2_1_wdata;
      end else begin
        ram_w32_l128_id2_1_rdata_out <= mem[ram_w32_l128_id2_1_addr];
      end
    end 
  end


endmodule



module madd_0
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_0
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_0
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_1
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_1
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_1
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_2
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_2
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_2
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_3
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_3
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_3
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_4
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_4
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_4
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_5
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_5
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_5
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_6
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_6
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_6
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_7
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_7
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_7
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_8
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_8
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_8
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module multiplier_0
(
  input CLK,
  input update,
  input [64-1:0] a,
  input [16-1:0] b,
  output [80-1:0] c
);


  multiplier_core_0
  mult
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c)
  );


endmodule



module multiplier_core_0
(
  input CLK,
  input update,
  input [64-1:0] a,
  input [16-1:0] b,
  output [80-1:0] c
);

  reg signed [64-1:0] _a;
  reg signed [16-1:0] _b;
  wire signed [80-1:0] _mul;
  reg signed [80-1:0] _pipe_mul0;
  reg signed [80-1:0] _pipe_mul1;
  assign _mul = _a * _b;
  assign c = _pipe_mul1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _pipe_mul0 <= _mul;
      _pipe_mul1 <= _pipe_mul0;
    end 
  end


endmodule



module multiplier_1
(
  input CLK,
  input update,
  input [64-1:0] a,
  input [16-1:0] b,
  output [80-1:0] c
);


  multiplier_core_1
  mult
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c)
  );


endmodule



module multiplier_core_1
(
  input CLK,
  input update,
  input [64-1:0] a,
  input [16-1:0] b,
  output [80-1:0] c
);

  reg signed [64-1:0] _a;
  reg signed [16-1:0] _b;
  wire signed [80-1:0] _mul;
  reg signed [80-1:0] _pipe_mul0;
  reg signed [80-1:0] _pipe_mul1;
  assign _mul = _a * _b;
  assign c = _pipe_mul1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _pipe_mul0 <= _mul;
      _pipe_mul1 <= _pipe_mul0;
    end 
  end


endmodule

